// ================================================================
//  Test-bench :  tb_modSwitch_qBBa_to_BBa
//                • ONE deterministic test only
//                • Uses the user-supplied stimulus / answer
// ================================================================
`timescale 1ns/1ps
`include "types.svh"

module tb_modSwitch_qBBa_to_BBa;
// ----------------------------------------------------------------
//  DUT I/O
// ----------------------------------------------------------------
logic clk = 0;
logic reset = 0;
logic in_valid;
logic out_valid;

rns_residue_t input_RNSpoly  [`N_SLOTS][`qBBa_BASIS_LEN];   // 22 residues
rns_residue_t output_RNSpoly [`N_SLOTS][`BBa_BASIS_LEN];    // 11 residues

// 11 (q)  + 11 (BBa)  = 22
localparam int QLEN   = `q_BASIS_LEN;        // 11
localparam int BBALEN = `BBa_BASIS_LEN;      // 11
localparam int TOTLEN = `qBBa_BASIS_LEN;     // 22

// ----------------------------------------------------------------
//  CLOCK
// ----------------------------------------------------------------
always #5 clk = ~clk;

// ----------------------------------------------------------------
//  DUT
// ----------------------------------------------------------------
modSwitch_qBBa_to_BBa DUT (
    .clk            (clk),
    .reset          (reset),
    .in_valid       (in_valid),
    .input_RNSpoly  (input_RNSpoly),
    .out_valid      (out_valid),
    .output_RNSpoly (output_RNSpoly)
);

// ----------------------------------------------------------------
//  USER–SUPPLIED TEST VECTORS  (constants)
// ----------------------------------------------------------------
localparam int NUM_TRIALS = 1;    // << only one run >>

// ----------  known input : 64 × 11  ---------------------------------
const rns_residue_t KNOWN_IN [`N_SLOTS][22] = '{
    '{0, 1139959117, 726617123, 939866751, 1101054909, 1910787954, 1082722200, 1953622552, 998113298, 876450072, 1661728428, 2112625357, 1419811165, 896997367, 1616153771, 1466324504, 1785119983, 2144932343, 943190406, 258722359, 1436875141, 1296049546},
    '{0, 1335435403, 776049247, 970384633, 965580893, 2095278784, 207766096, 392990415, 2013836012, 705465416, 107591171, 218718128, 715799810, 46960383, 372403674, 101379032, 206989336, 741514970, 1864878476, 1874591947, 1565085699, 705825841},
    '{0, 1009092702, 645052409, 727448244, 1392135697, 324874751, 1287008776, 885210078, 760099671, 1347830250, 2128704505, 1803290161, 1557017431, 604579136, 1167265685, 20017128, 1578375818, 1809351894, 362698446, 255849229, 1892899298, 757278422},
    '{0, 1834084134, 2120337403, 2013836257, 103324888, 1134380307, 1605367068, 274292550, 1890007266, 884872490, 2137966810, 1196363765, 1416180165, 329578282, 2101893320, 294500171, 1968395373, 70754716, 1116754073, 476509903, 1416017618, 1822388973},
    '{0, 379133673, 1091876763, 1286543723, 999529156, 198306960, 1037441904, 56853492, 1767465038, 320821531, 1573856523, 1658840261, 395652189, 1931625719, 1855753628, 2054141357, 560767632, 1521592835, 886379865, 201884305, 2030906232, 299912295},
    '{0, 1338185242, 1228946350, 34865958, 1988573395, 141063649, 1024934630, 2072113756, 484022250, 134639499, 1596277839, 2137406913, 330282610, 294222474, 461442131, 308338653, 2070408484, 1938542747, 736685720, 2004200242, 2087574198, 995944841},
    '{0, 33294222, 775717376, 589871314, 182377984, 912476422, 807722535, 401137798, 1132037772, 1847691905, 809159092, 1715971898, 1843997340, 2010042794, 721516478, 1964728612, 1616343162, 1106270932, 525588396, 1806909312, 1534017930, 752060495},
    '{0, 822108697, 300935668, 1840383577, 1992678590, 1966625411, 488731659, 1316442019, 2041909422, 1826676692, 1379496565, 920690674, 65507198, 131204130, 310740154, 228785546, 216783516, 1407727966, 714786077, 857072597, 34276179, 984072861},
    '{0, 930669969, 170594468, 1700853867, 286544209, 1197491185, 1253233675, 866391137, 350135641, 1484233798, 1277651821, 85622950, 193306148, 1830705940, 901768701, 1991480198, 1219816283, 426933459, 99027926, 1721535947, 1733644898, 527857612},
    '{0, 1811838908, 1896834477, 1366575519, 2002428613, 1159918619, 1657340327, 1513257506, 1338887090, 1589867022, 1816564077, 750797806, 182244896, 841420117, 1116438639, 2021539257, 1308886423, 656722289, 1666813904, 1751424712, 1645276986, 181079512},
    '{0, 415895252, 1057916259, 875519619, 1852423673, 197512480, 1509359114, 952229989, 1747062584, 1585099667, 1459258917, 1222413081, 199665866, 1248064040, 680876413, 1699691383, 1907037542, 1111947112, 1731731250, 1316636595, 1949002514, 1809002182},
    '{0, 1807632617, 1195838340, 980159495, 2054775305, 855678120, 1074190186, 1880788757, 1862727606, 856074675, 81790953, 1242586049, 850384948, 870986249, 439959291, 184374327, 1627286655, 1088284440, 152223217, 780288244, 1013035417, 496780647},
    '{0, 267090854, 1433431741, 688452547, 342651797, 527468934, 1766984766, 1986737785, 188941817, 852584550, 1279267193, 206116495, 1346636882, 526283129, 1493045004, 207395922, 921178065, 1010016110, 1568328287, 1673743485, 477635592, 1818243596},
    '{0, 998749039, 1322844086, 881652989, 308233099, 1865664012, 609634034, 1291270222, 1173647682, 1508991253, 317136011, 651907553, 786362613, 988886266, 1434526243, 1801964092, 1762412562, 1992350648, 2099829554, 1437068038, 253953529, 879636361},
    '{0, 560984648, 1387647553, 1953927620, 624312929, 1580864956, 106261725, 614736243, 944575835, 889837992, 1414038366, 233948629, 2143824226, 2016465607, 433589157, 700504935, 1256423303, 1232495516, 242356673, 38884406, 1770992584, 1392499332},
    '{0, 696393614, 2117283842, 1734667903, 675230518, 787070613, 776120282, 950474387, 1938616435, 1824902343, 604167412, 238789046, 1806764561, 1402045716, 533739188, 218676578, 1513966179, 1731134314, 443528406, 1707018194, 1845812234, 883222725},
    '{0, 566086066, 2075192066, 1638895466, 1019700008, 1249469817, 653177944, 1690230537, 136180606, 1864732447, 579508602, 1350497354, 2099121824, 1896473863, 480080596, 767401629, 1524547031, 1127372772, 885857549, 1617756519, 1525540109, 671755927},
    '{0, 767856670, 673328982, 1191367268, 636775229, 163111809, 1799502421, 2119291510, 749963837, 72983111, 463032457, 1609799384, 26430894, 1122956748, 1356873884, 110005457, 59982106, 688808259, 354904861, 1701293100, 1291485073, 1743982977},
    '{0, 506462505, 979378226, 1587813312, 1122504690, 466124310, 106352777, 518076220, 1879256982, 1774722806, 375234760, 41597010, 1454984900, 815254894, 185209172, 1651373626, 1877895155, 67697567, 1525210764, 1931618465, 1550824021, 1919926544},
    '{0, 1240000159, 172773677, 1440542585, 1930438077, 1088835941, 702024211, 520986392, 1890842376, 1013303489, 128361299, 132581080, 1713441843, 674096212, 1783145875, 1041125556, 1015255268, 1288048784, 562855182, 556979282, 188047061, 1213226792},
    '{0, 275672181, 1872825888, 515444028, 1089438314, 874494124, 543391690, 579414763, 1474932108, 41695289, 998643963, 1199642453, 933605252, 620126902, 1328314659, 954971329, 603313924, 1235842627, 2078452120, 1618169082, 2075036318, 1916785840},
    '{0, 99404516, 1289920812, 886474194, 1149666510, 243098004, 1143177077, 1502624603, 1326790141, 942202483, 2015643760, 357873327, 1671149772, 1964582802, 20485058, 741334218, 2048140651, 1369076848, 1292710338, 749684792, 555477529, 1093387084},
    '{0, 2049751032, 1155836750, 354964871, 1641244976, 1831229493, 779841756, 1674478295, 45674298, 1174910631, 325174890, 1729773150, 2023869336, 1090875361, 1074889835, 268901298, 1565350926, 1808428014, 755995804, 432443514, 566881430, 1107640352},
    '{0, 918967290, 1634854097, 943766488, 2071106284, 1059779381, 1471096060, 867279598, 1064347435, 1410785241, 1292626625, 1152780468, 1090143291, 1045337198, 57013159, 788443168, 692151279, 1051879514, 936772660, 1292398236, 357477852, 604469681},
    '{0, 1073688997, 1444168241, 1099494586, 17802383, 566369860, 1696723703, 1416322135, 1424427914, 260552178, 927591220, 533917909, 25758009, 922840270, 657474210, 1267606443, 525738659, 1642950338, 1807232156, 1759482028, 1599869973, 894549898},
    '{0, 712920507, 1166971371, 1070221267, 988930622, 1533589943, 268994942, 1467673016, 743651510, 299349664, 1261366936, 201249629, 842042696, 463353426, 239953777, 2000461156, 1198192560, 533447611, 855098220, 1210110081, 689294022, 496517864},
    '{0, 818138195, 241180357, 1297256065, 1417398954, 208215361, 1152960505, 788267793, 1269713765, 1568957478, 1175362919, 1315203289, 943146550, 977570704, 387746458, 1764343842, 290252053, 434541080, 286378600, 1811547599, 1905687658, 1582393337},
    '{0, 1209336991, 1310345311, 1536311626, 476650948, 1121733160, 722236522, 1369852357, 641287507, 810244105, 658686053, 401812781, 433724346, 480564376, 1674703786, 925445394, 935296222, 327194589, 1298550041, 666778106, 1325241718, 76643607},
    '{0, 657049995, 1091564320, 752944434, 1920698776, 357895561, 1085348981, 1557806845, 1794051942, 1089796782, 2073975964, 367746363, 1928545634, 1015105149, 1600526927, 354631055, 1418256911, 1073252103, 726926993, 1896206873, 1572737305, 1324205866},
    '{0, 1962775112, 1899908485, 1836559178, 935481040, 1717773706, 203309299, 1821963343, 1363313735, 427436306, 1393168694, 772611700, 783666504, 1356658985, 1346315000, 1376036285, 387769097, 230666972, 1424190621, 1686793981, 1998690901, 1348803997},
    '{0, 113119730, 1003221961, 1249049316, 9104725, 1092212996, 757168158, 1149165080, 817687436, 847214826, 898650606, 439293021, 1333992651, 1348594590, 1378183215, 997327964, 1979496535, 1038350652, 1215046943, 1645664326, 1885945995, 1998069001},
    '{0, 541813567, 96059842, 1816140693, 1199077579, 517973403, 1549472049, 283257220, 250627822, 1688027794, 655393001, 1634038068, 1555185189, 568938406, 2122106802, 225408848, 61555520, 1377515087, 1174468927, 985343669, 1516254778, 748302916},
    '{0, 443706352, 1305089481, 1382576642, 1814558850, 970632717, 77620500, 1849647958, 166746383, 189646627, 1713465405, 449015366, 1453258100, 766514869, 812998044, 2124639178, 726199487, 33849921, 892037025, 925398373, 1645003507, 639565206},
    '{0, 1353583770, 737236629, 1564380070, 2081434930, 1231938720, 1287087218, 1529542961, 1505435945, 274506470, 1390014222, 1461034080, 1145232095, 1335470782, 1715392967, 673879267, 365210216, 995567478, 1374775367, 1533219402, 2062280973, 246421527},
    '{0, 1583834681, 13990921, 596510581, 101157579, 1819326018, 626777152, 1710485859, 384573419, 1660090007, 1366134627, 115915885, 1419937466, 435385132, 469181677, 595107849, 77876203, 2011442759, 1160319160, 1178062700, 624789641, 1035187175},
    '{0, 519295113, 38506597, 713944731, 1912725123, 689678170, 2092575163, 621425520, 1143681514, 1098368957, 2145791686, 558867749, 567666957, 479838541, 197126848, 107021419, 474736717, 197974097, 393294548, 441265304, 1036961893, 395324699},
    '{0, 1762187035, 594753672, 289760556, 1293552920, 970563251, 1723335556, 134635611, 1675706945, 1552190255, 483091807, 1975977725, 223178470, 1174040890, 1118595292, 1952444345, 1826079565, 605898426, 1301921145, 835906286, 1541134747, 1474331085},
    '{0, 2114815633, 2013395761, 1449436477, 1132328872, 70509075, 241240563, 2113659245, 1221886035, 329111807, 95253013, 294127811, 62162323, 495959732, 1902740243, 1233464688, 467733513, 109515319, 1633646835, 1024579210, 1134994380, 1817411694},
    '{0, 1189227031, 1769725161, 1145925244, 212015362, 1216551449, 1641017464, 701407668, 1136213647, 114993386, 460079681, 1296952185, 1351527828, 1590696031, 1773741044, 1308579672, 574041636, 1086895747, 995786407, 2062439827, 1579966796, 2123642340},
    '{0, 1879082276, 332408959, 1145383539, 1678737552, 1363654152, 1775975936, 945449474, 1239516572, 2087772428, 668157536, 2095960587, 79033491, 1428144688, 1438338376, 2142779985, 865300978, 1240196310, 264138255, 1593426634, 543065275, 225493889},
    '{0, 1178700778, 1133490373, 1911650388, 453590396, 331099592, 791184821, 40119829, 651916464, 990806038, 1812981207, 1095221814, 1190586311, 438172465, 1477583327, 1693298016, 146593409, 1793117245, 1138146960, 2059309070, 1179204489, 421254160},
    '{0, 1457460237, 550124273, 231540297, 2146263398, 57371577, 368706914, 731891440, 1241331803, 251069418, 1590943970, 2023962815, 769002186, 656272126, 1609893051, 6981110, 16680821, 1463920769, 2058299732, 1651530526, 1463690146, 1283706803},
    '{0, 1226309268, 1649608779, 1452190276, 500560720, 1707877178, 1973769689, 1590816965, 701465182, 223432210, 1146292910, 106133788, 1413943752, 1826925851, 339311634, 894489849, 1341563554, 2009226640, 1997060509, 1253022896, 1131472573, 1134547736},
    '{0, 197047463, 1988751714, 2198910, 385198704, 686955728, 530178958, 1838788453, 94212402, 406553955, 556678523, 1240623188, 1686732973, 1535332682, 1889979129, 823302541, 116531031, 1694477324, 1229944355, 439567622, 2082087753, 1759278908},
    '{0, 1075690737, 1733936180, 246255412, 84046831, 562804286, 1969456709, 654282535, 431387402, 775579303, 1402399369, 1823468170, 2109496064, 588973622, 20660936, 707135981, 1215664934, 1668584035, 890231140, 409790666, 1606906814, 1860208185},
    '{0, 482167408, 749199826, 223931436, 211607537, 598537986, 1463595174, 825271886, 1720693193, 1952927478, 1358335396, 412444327, 1974082437, 34601887, 138932163, 402979255, 1446297925, 1398043725, 1179283040, 1939343553, 796258527, 779325374},
    '{0, 1368710193, 1010223426, 832945983, 1904089518, 1256107533, 1126383548, 1573381021, 338980883, 1793851485, 1411010571, 1942132626, 90963370, 1110449145, 1907683657, 1399254405, 1361923948, 315420873, 36432409, 1354611674, 261340385, 725945562},
    '{0, 1711391996, 1832373192, 1400186781, 2069604702, 445619896, 1937725586, 317734786, 628543401, 1654142290, 2049370848, 778421544, 902292472, 807349210, 784438419, 2140171397, 781689787, 1668371710, 1816416933, 2025830740, 549112336, 1091561311},
    '{0, 2001363630, 1569584639, 2738540, 1406402323, 1875249127, 1884751605, 813875558, 416104000, 1223520321, 407466589, 1133723932, 2056823668, 591163356, 1798821345, 1351176593, 1738855035, 1438121748, 1302177609, 2045558694, 1252622574, 1320529914},
    '{0, 944131141, 1679881521, 137078133, 218169602, 499650478, 1427968864, 545133608, 2128283499, 1751463290, 1505090877, 378336277, 1805836639, 1201833262, 482858671, 1199831630, 221166162, 1517777793, 282587605, 1415180062, 649731308, 288593939},
    '{0, 2141701456, 889447512, 595275329, 1757164137, 1767467753, 1084794503, 1945688084, 725652453, 1840046374, 2139500253, 180882270, 2111355394, 2086666344, 1120058663, 1944068699, 1244533602, 391341901, 617724405, 376800875, 428265513, 278303433},
    '{0, 1841460212, 408268047, 44849044, 986446520, 830522490, 1215996098, 1944728640, 1092612267, 1345630060, 1240636009, 2143855708, 1180131442, 1015372460, 2130461058, 667867688, 142102080, 743637836, 47728946, 236574515, 152320764, 98317257},
    '{0, 1916526861, 2032945812, 158471968, 478363369, 1347634242, 116637503, 1982033075, 517039521, 2064659788, 1114216459, 2111626738, 590350442, 2095434731, 395508774, 273215865, 553999621, 204908461, 905875390, 1007398326, 163193034, 122128591},
    '{0, 599287523, 2048032231, 119480112, 1207892124, 1365397780, 1791430912, 1399718973, 317074422, 1390923349, 129186018, 830105334, 2140043092, 484200085, 16548072, 2080540313, 1053378684, 1514496024, 940696051, 1503615405, 2116595367, 56843714},
    '{0, 1453208562, 2022047013, 1756129893, 357250158, 361144691, 1694834217, 1972344402, 2127382757, 208073152, 995348361, 950953474, 61601199, 795035125, 1801725367, 610372563, 1438572094, 1908959765, 1663738360, 709873932, 1038185067, 578292259},
    '{0, 768268797, 672058135, 48860939, 1350791639, 370977499, 1706052991, 1341134442, 1658726665, 2079434427, 1419314168, 1969524065, 977286439, 1901656550, 1121195610, 560976971, 1522582203, 861521188, 537027713, 1461794069, 2014770649, 1512363050},
    '{0, 281885187, 666650009, 1482637256, 725412614, 426349625, 649900130, 1518113779, 1508540972, 239299258, 444107125, 103228968, 139468394, 1401679318, 1296984322, 2138359612, 1935447756, 1511103412, 318970920, 2134640065, 1090281154, 1794683575},
    '{0, 1023187644, 513626984, 1583018684, 1359535150, 2077302849, 1970755429, 104708138, 1169222227, 2023740551, 1044336559, 2029621937, 1120253955, 1302634413, 376909947, 1057593122, 110318203, 686648303, 1955322227, 1820319609, 1594848230, 352437225},
    '{0, 1000217728, 1359042055, 710906063, 2039936923, 999758695, 1928316656, 2050383286, 1227345332, 2567439, 1958758582, 102666544, 825339635, 1941562881, 2039557320, 2015581026, 2017493768, 769497420, 1091187933, 626877467, 1062073927, 1347258552},
    '{0, 1861084514, 1713882088, 1450070099, 460951795, 1824103046, 859760768, 275519517, 1719398220, 965264600, 800754342, 1682990973, 2133449586, 1681766549, 1291392480, 1672480744, 1421287134, 1069072489, 243339522, 334791914, 1632990877, 1656507348},
    '{0, 920539188, 179146124, 1409150951, 920089857, 1657283740, 889662516, 2122931353, 1441715982, 1573423885, 1843703831, 388808798, 987845365, 167663574, 2067765902, 1984540332, 686758178, 846343994, 1533898167, 1572325057, 511498072, 679811224},
    '{0, 1821191953, 1322208162, 162979028, 1127620014, 547610980, 773418938, 1136412453, 654561708, 835414208, 644693037, 1267694532, 1914384905, 357870488, 1899565469, 1667705793, 1553932041, 2113082891, 329890217, 2131566736, 1036101988, 490438852},
    '{0, 1596542719, 337228497, 1714592618, 1342318162, 1094140098, 728754077, 1025726344, 807611204, 2065238405, 929712599, 402409253, 220587165, 443285300, 1823477731, 1047125085, 557292329, 633481815, 1730201201, 1264859085, 746459006, 1264664728},
    '{0, 2046676616, 1930345071, 2047193936, 2123866676, 409673837, 1043454822, 2006228434, 290591003, 824732323, 1218388965, 2116775999, 520455172, 786533712, 1411999376, 377274974, 487230736, 1526590878, 906545918, 405178767, 1681392247, 208102737}
};

const rns_residue_t KNOWN_OUT [`N_SLOTS][11] = '{
    '{2406575, 313906966, 605474624, 934239537, 1589668363, 1567356734, 1471776138, 364225185, 1613769651, 1153893135, 1856411822},
    '{81001096, 511913739, 1130195616, 935905454, 1510787025, 1859042182, 520698806, 141283181, 957394802, 1041317308, 273885315},
    '{2055992580, 1531891891, 1090933461, 572525100, 1245624002, 287953027, 1925629873, 1565019550, 1660605871, 516066792, 1970769398},
    '{680468203, 1402207188, 847597246, 956089897, 1994455403, 402658697, 1729960384, 1444148079, 1247481335, 104546859, 911579519},
    '{1981331186, 270691168, 578111836, 1485776934, 523322228, 1672899391, 581071596, 209906933, 1937820572, 1722258337, 656554988},
    '{1507789192, 1057874066, 1239533268, 1520038621, 618026960, 637922026, 366521069, 1066877968, 154029783, 266603930, 1749384995},
    '{939961214, 1362239244, 258100131, 635551601, 33265343, 1987051861, 1182272113, 963446960, 1728519845, 592150413, 1185632388},
    '{1459793209, 1114861983, 1708067667, 233711142, 1053016725, 1253721065, 1355798783, 45355269, 708739769, 130643320, 396704188},
    '{1235861497, 1141593479, 1040232804, 1310947662, 1551004462, 744998938, 655539971, 802686368, 326224097, 1070548522, 315525028},
    '{719126444, 1986038605, 1624781605, 1205748015, 578864915, 792759487, 1887702220, 1954252474, 842445442, 2041960974, 1171648770},
    '{993668077, 1208123452, 1870638289, 1437634358, 1217623833, 1817907176, 364254771, 2034380733, 1861736132, 1836298811, 1008315771},
    '{531244676, 176969436, 499291796, 919046049, 363811625, 1243783645, 2093180313, 113600263, 1858652316, 1521120752, 766368520},
    '{512137188, 262417205, 753660508, 996624964, 1438329733, 1707058579, 1561088649, 1973453196, 1026946607, 1195063626, 897700266},
    '{1492782280, 1877260613, 725974715, 2114713929, 1886993401, 1006122773, 64064158, 4562261, 389883655, 1452813470, 140368152},
    '{973137646, 448824411, 1273111477, 1073719071, 124623805, 222994203, 676132011, 147163343, 983114351, 1168296970, 1424746320},
    '{1760891879, 489222995, 1161239651, 611599488, 1369000515, 1880566775, 407302070, 1765713593, 1850035282, 1671526585, 650239463},
    '{99592340, 402659615, 1136250757, 153344595, 539961838, 1017773168, 1351528001, 1903210076, 1127800961, 942725257, 2144914371},
    '{356720379, 726306145, 841674202, 1513398140, 1675121933, 2051788094, 1636822034, 1504253498, 677505606, 1726797323, 431762233},
    '{1797078652, 965189296, 2101889306, 2036607256, 1629679618, 1516407549, 647705664, 141529315, 343187844, 1134852132, 793334257},
    '{1697693148, 602810806, 347465435, 585980505, 957143300, 618156830, 727220297, 1091530320, 90661765, 1315135908, 1392059309},
    '{54406186, 1641040526, 172420453, 20348990, 658270238, 380429789, 767586555, 1925354464, 982583157, 783985997, 782395249},
    '{1360751317, 1221793502, 1655693209, 2032112247, 199413, 1102406212, 2074409899, 1391658613, 1232458906, 1413409323, 1984506769},
    '{1015913994, 194203877, 996827189, 1295829275, 2142890934, 1609431404, 1662833724, 24006374, 1029637171, 1162709024, 1076173463},
    '{414133899, 1054077184, 1522311628, 1266050552, 340419067, 92322600, 1952973300, 769560695, 1233956586, 696948476, 1665236991},
    '{1905660568, 108391766, 686072115, 1169578648, 1369767692, 479475575, 1276715384, 1639168422, 197997224, 2122651339, 2106704340},
    '{2146204958, 1893340932, 2033795022, 854911643, 600729427, 1915012376, 475674864, 1944663921, 158512527, 1748072582, 1858882740},
    '{1256330565, 1363158609, 550996612, 965644187, 655911434, 1442701579, 397793942, 804160830, 2023525790, 1485967739, 1986138205},
    '{790536360, 576932890, 408926549, 608054726, 1037418890, 1035668867, 473407492, 1999421932, 402191142, 64965890, 2017865625},
    '{1066811454, 487286723, 1473468771, 91359911, 1741399031, 2091868701, 1989685199, 834080369, 1295874215, 867456099, 1689179528},
    '{1095444225, 1689395509, 454423238, 756358769, 1761802148, 1556338264, 256421482, 752261882, 1563366245, 587761475, 329435887},
    '{704614972, 628351179, 2123456575, 689287272, 1413576382, 1256201973, 1575448078, 413991834, 579738227, 690582911, 1788497851},
    '{1263759218, 1224427145, 497561573, 2041789324, 525661179, 37790758, 1074328797, 1471993313, 1289280764, 1781870380, 1674283996},
    '{734086029, 1496252073, 1545358428, 517601706, 590606257, 1582342532, 2068120328, 169232049, 1451417623, 1918733375, 169362086},
    '{440875221, 211096, 1975290762, 1864165673, 2132420018, 1997881216, 207978271, 297358748, 223630192, 1296401166, 1132842309},
    '{690969991, 425860733, 613422242, 1169018016, 631200332, 1628298016, 471598227, 1590758801, 1642195566, 71755622, 1598666286},
    '{1064509008, 1171851795, 1664557051, 944936064, 532990375, 1362573797, 1041741186, 1822302322, 1031694695, 907367624, 541551278},
    '{399265170, 644856550, 774293876, 1156413635, 1832643562, 66869645, 1810055000, 705985050, 922869234, 482276845, 198385014},
    '{1597192379, 1793492906, 394564745, 1567243632, 1661645748, 854528972, 1307780663, 1171051708, 1279202903, 939443532, 1519436909},
    '{1287479889, 592383651, 757140919, 986077766, 197728418, 1496347989, 1076023385, 310639074, 1944694510, 1841349452, 1781596949},
    '{877293530, 680735415, 1276096439, 1320432424, 682780658, 245032395, 364988159, 393689510, 1414584694, 106383080, 212476702},
    '{76890534, 1463999637, 1682399220, 312822740, 700779533, 1066818239, 1049517706, 1615351145, 1685240303, 335888525, 2080584363},
    '{1276474204, 281092366, 882130565, 1646368213, 1079802398, 530530517, 218465760, 1825414618, 1328024520, 596714516, 1589355981},
    '{1904784871, 2018720024, 826138003, 897162357, 296692050, 624870, 1522206850, 1573945787, 942611545, 699724978, 1480432030},
    '{172168037, 956953317, 1141769605, 124628910, 81326518, 1744788010, 176857354, 702079915, 1192436350, 1420610320, 1013178392},
    '{795428645, 165369361, 1413723967, 317211378, 126869386, 2139089952, 1910725768, 1183584878, 951374247, 212440062, 991754962},
    '{550123113, 1176413791, 943939508, 944683965, 1098339517, 1155793733, 29380478, 1292246679, 1359073312, 1420581464, 115591543},
    '{1097670016, 920110368, 992106981, 392351802, 1741179579, 1504664780, 1083176042, 1607075061, 72701877, 490662662, 375538199},
    '{853297895, 1549249585, 676457627, 1848545344, 386240396, 709855208, 1066061302, 540213286, 2048147107, 1956987137, 927762976},
    '{1323850257, 164774676, 1678604188, 1953881943, 2062196185, 589043076, 1984699685, 524787334, 1956415317, 917888968, 225000876},
    '{727123941, 1010281021, 1547777933, 882506301, 831072733, 103561200, 1934965260, 2096307526, 682153045, 790133528, 1296402548},
    '{1189060403, 998859921, 1777087363, 1599721371, 1517257180, 1791045272, 187718463, 529070739, 1367756034, 735762285, 1164915924},
    '{1642288113, 2149147, 1194360260, 1593755617, 1287594959, 1327956309, 2142396084, 1142970209, 1468627592, 1166401127, 1005490367},
    '{1883487776, 1721982432, 1449901647, 35967890, 167599815, 2042122320, 1994596462, 1576198708, 808116175, 494991200, 1327915565},
    '{1737756517, 75181361, 250878390, 330465822, 2025578758, 1376875783, 388786945, 1658435564, 1633453352, 304563362, 792004994},
    '{1121753646, 1955676666, 2091500489, 236897374, 394681111, 778270610, 1698553150, 1962482671, 506902708, 714000722, 1942692519},
    '{1046961526, 1032807288, 1201942487, 1456638309, 48840388, 372821246, 686716535, 55738262, 2059014790, 1649686815, 431303318},
    '{856024551, 1126229164, 1158287201, 1340354664, 1493953049, 933558923, 1331379471, 1843382751, 2064308379, 2010055463, 1884754857},
    '{569350354, 338377234, 902771092, 267012725, 912847616, 1341904049, 1742999534, 791530456, 266951401, 23151614, 780811672},
    '{445401295, 698297736, 22414416, 1537993602, 731951509, 212997683, 1649163198, 1338983511, 6556059, 609123505, 1419375288},
    '{454542236, 1841160733, 1625951161, 106803849, 1207382414, 1346454852, 1769967665, 1285718905, 60631945, 1661393899, 994437922},
    '{666346933, 489194288, 879451083, 709680126, 2144914019, 1470930075, 1604786121, 1706382111, 1524219264, 1988380883, 1002808500},
    '{1171553528, 1012450913, 438759822, 976368811, 1731737561, 1750967259, 301582012, 1659309318, 1091393147, 60892554, 984982174},
    '{1495411137, 1638380283, 866160050, 790454697, 1753231758, 960718445, 1928281240, 1972799288, 1951001614, 1453127537, 966844749},
    '{1737016703, 598355960, 606607430, 388968163, 1080018074, 238100719, 36803152, 1026589462, 1393076867, 698860141, 1205040083}
};

// ----------------------------------------------------------------
//  TEST PROGRAM
// ----------------------------------------------------------------
rns_residue_t golden_answer [`N_SLOTS][`BBa_BASIS_LEN];
bit          mismatch;
int unsigned pass_cnt = 0;
int unsigned fail_cnt = 0;
logic DEBUG_MODE = 0;
initial begin
   // ----------- reset ------------
   @(posedge clk);
   @(negedge clk);
   reset    = 1'b1;
   in_valid = 1'b0;
   @(negedge clk);
   reset    = 1'b0;

   // *************************************************************
   //  ONLY ONE TRIAL – load the static vectors
   // *************************************************************
   for (int k = 0; k < `N_SLOTS; k++) begin
      // copy q-part
      for (int j = 0; j < QLEN; j++) begin
         input_RNSpoly[k][j]        = KNOWN_IN [k][j];   // q residues
         input_RNSpoly[k][j+QLEN]   = KNOWN_IN [k][j+QLEN];   // BBa residues (kept)
         golden_answer  [k][j]      = KNOWN_OUT[k][j];   // expected BBa result
      end
   end

   $display("\n\n");
   if(DEBUG_MODE) begin
        //$monitor("to_be_dropped_RNSpoly 0 1 = %0d", DUT.to_be_dropped_RNSpoly[0][1]);
        //$monitor("xhat_f 0 0 =%0d | " , DUT.xhatf_fastBconv_output_RNSpoly[0][0]);
        //$monitor("xhat_f 0 1 =%0d | " , DUT.xhatf_fastBconv_output_RNSpoly[0][1]);
        //$monitor("xhat_f 0 1 =%0d | " , DUT.xhatf_fastBconv_output_RNSpoly[0][1]);
        $display("input 0 0=%0d, input 0 11 =%0d | " , DUT.input_RNSpoly[0][0], DUT.input_RNSpoly[0][11]);
        $display("drop 0 0=%0d, drop 0 1 =%0d | " , DUT.to_be_dropped_RNSpoly[0][0], DUT.to_be_dropped_RNSpoly[0][1]);
        $display("chi 0 0=%0d, chi 0 1 =%0d | " , DUT.to_be_kept_RNSpoly[0][0], DUT.to_be_kept_RNSpoly[0][1]);
    end

   // -------------- Drive DUT -----------------
   @(negedge clk);
   in_valid = 1'b1;
   @(negedge clk);
   in_valid = 1'b0;

   // -------------- Wait for result -----------
   while (!out_valid) begin
      @(posedge clk);
   end
   @(posedge clk);

   // -------------- Compare -------------------
   mismatch = 0;
   for (int k = 0; k < `N_SLOTS; k++) begin
      for (int j = 0; j < BBALEN; j++) begin
         if (output_RNSpoly[k][j] !== golden_answer[k][j]) begin
            //$display("[%0t]  SLOT %0d  RES %0d  MISMATCH  DUT=%0d  GOLD=%0d", $time, k, j, output_RNSpoly[k][j], golden_answer[k][j]);
            mismatch = 1;
         end
      end
   end

   if (mismatch) fail_cnt++; else pass_cnt++;

   // -------------- Summary -------------------
   $display("\n==================================================");
   $display("Mod-Switch deterministic test finished");
   $display("      Passed : %0d", pass_cnt);
   $display("      Failed : %0d", fail_cnt);
   $display("==================================================\n");
   $finish;
end

endmodule