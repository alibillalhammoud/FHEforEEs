`ifndef TYPES_SVH
`define TYPES_SVH

// ---------------------------
// Basic data types
// ---------------------------



// NTT
`define BASE      32'd2
// Width of each RNS residue (one small prime)
`define RNS_PRIME_BITS 32
// RNS residues
typedef logic [`RNS_PRIME_BITS-1:0] rns_residue_t; 
typedef logic [(2*`RNS_PRIME_BITS)-1:0] wide_rns_residue_t;
// Vector / slot params
`define N_SLOTS   64
// moduli and RNS bases
`define t_MODULUS 257

`define q_BASIS_LEN 11
//`define q_MODULUS = 536092687689737712660299305370020840707037344303743567681198293980556215074372863278673727266177
parameter rns_residue_t q_BASIS [`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353};
//`define B_MODULUS = 2086045702160390514072457421164142647843268814746900546792219301529141418454085790414389880321
`define B_BASIS_LEN 10
parameter rns_residue_t B_BASIS [`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337};
//`define Ba_MODULUS = 2147503489
`define Ba_BASIS_LEN 1
parameter rns_residue_t Ba_BASIS [`Ba_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147503489};
`define qBBa_BASIS_LEN 22
//`define qBBa_MODULUS = 2401582888476023779443294070753805757615044045174800139284098902756577490274881128570727198734820745298450301532339857214864378319647024214690248526201090429246246041638715397173165827069546764128513
parameter rns_residue_t qBBa_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353, `RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147503489};

// RNS integers
typedef rns_residue_t rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef rns_residue_t rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef rns_residue_t rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
/*typedef rns_residue_t rns_coef_qBBa_BASIS_t [`q_BASIS_LEN + `B_BASIS_LEN + `Ba_BASIS_LEN];*/
// Polynomials
typedef rns_int_q_BASIS_t q_BASIS_poly [`N_SLOTS];
typedef rns_int_B_BASIS_t B_BASIS_poly [`N_SLOTS];
typedef rns_int_Ba_BASIS_t Ba_BASIS_poly [`N_SLOTS];
/*typedef rns_coef_qBBA_BASIS_t qBBa_BASIS_poly [`N_SLOTS];*/
// wide RNS integers (each residue is double the length for mult)
typedef wide_rns_residue_t wide_rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
// wide Polynomials
typedef wide_rns_int_q_BASIS_t wide_q_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_B_BASIS_t wide_B_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_Ba_BASIS_t wide_Ba_BASIS_poly [`N_SLOTS];

// ---------------------------
// precalculated values
// ---------------------------
// Example constant “twist” factors (all 1s for now)
parameter rns_residue_t twist_factor   [`N_SLOTS] = '{default: '1};
parameter rns_residue_t untwist_factor [`N_SLOTS] = '{default: '1};

// fastBConv precalculated inverses
parameter rns_residue_t z_MOD_q[`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1340848717, `RNS_PRIME_BITS'd1950706637, `RNS_PRIME_BITS'd136505383, `RNS_PRIME_BITS'd1261863396, `RNS_PRIME_BITS'd490720514, `RNS_PRIME_BITS'd2048232271, `RNS_PRIME_BITS'd561180295, `RNS_PRIME_BITS'd2064343317, `RNS_PRIME_BITS'd1284162414, `RNS_PRIME_BITS'd426116969};
parameter rns_residue_t z_MOD_B[`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd400603566, `RNS_PRIME_BITS'd1317047788, `RNS_PRIME_BITS'd1877527982, `RNS_PRIME_BITS'd816591707, `RNS_PRIME_BITS'd1500256234, `RNS_PRIME_BITS'd8640588, `RNS_PRIME_BITS'd1509953789, `RNS_PRIME_BITS'd1256593971, `RNS_PRIME_BITS'd1660146682, `RNS_PRIME_BITS'd390117507};
parameter rns_residue_t y_q_TO_qBBa[`qBBa_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1514938357, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1663002026, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1202970911, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1254269319, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd15070697, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd93592423, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd345241794, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd126359634, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1571891470, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1004678308 },
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};
parameter rns_residue_t y_B_TO_Ba[`Ba_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd33728781, `RNS_PRIME_BITS'd1756228743, `RNS_PRIME_BITS'd487215260, `RNS_PRIME_BITS'd501135696, `RNS_PRIME_BITS'd459470026, `RNS_PRIME_BITS'd1877657833, `RNS_PRIME_BITS'd50297305, `RNS_PRIME_BITS'd56214635, `RNS_PRIME_BITS'd1200871039, `RNS_PRIME_BITS'd1750218591 }
};
parameter rns_residue_t y_B_TO_q[`q_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd10, `RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd92 },
'{ `RNS_PRIME_BITS'd1219156511, `RNS_PRIME_BITS'd1608499681, `RNS_PRIME_BITS'd371154937, `RNS_PRIME_BITS'd924754142, `RNS_PRIME_BITS'd2003633539, `RNS_PRIME_BITS'd627440795, `RNS_PRIME_BITS'd1066486116, `RNS_PRIME_BITS'd1296251710, `RNS_PRIME_BITS'd1679092476, `RNS_PRIME_BITS'd772683368 },
'{ `RNS_PRIME_BITS'd1367502590, `RNS_PRIME_BITS'd1413619003, `RNS_PRIME_BITS'd1604587363, `RNS_PRIME_BITS'd796115568, `RNS_PRIME_BITS'd154115966, `RNS_PRIME_BITS'd287007179, `RNS_PRIME_BITS'd457558717, `RNS_PRIME_BITS'd43558045, `RNS_PRIME_BITS'd1825868505, `RNS_PRIME_BITS'd2117666329 },
'{ `RNS_PRIME_BITS'd488607457, `RNS_PRIME_BITS'd725589953, `RNS_PRIME_BITS'd166254356, `RNS_PRIME_BITS'd1679376923, `RNS_PRIME_BITS'd375851890, `RNS_PRIME_BITS'd962572449, `RNS_PRIME_BITS'd40302594, `RNS_PRIME_BITS'd37730088, `RNS_PRIME_BITS'd1726493613, `RNS_PRIME_BITS'd1162981935 },
'{ `RNS_PRIME_BITS'd317361695, `RNS_PRIME_BITS'd1920884754, `RNS_PRIME_BITS'd1303976625, `RNS_PRIME_BITS'd107931280, `RNS_PRIME_BITS'd1804980561, `RNS_PRIME_BITS'd1467513527, `RNS_PRIME_BITS'd1597511531, `RNS_PRIME_BITS'd1771541117, `RNS_PRIME_BITS'd2104139963, `RNS_PRIME_BITS'd695454200 },
'{ `RNS_PRIME_BITS'd875545508, `RNS_PRIME_BITS'd1106807570, `RNS_PRIME_BITS'd531200008, `RNS_PRIME_BITS'd656659131, `RNS_PRIME_BITS'd318605813, `RNS_PRIME_BITS'd571007940, `RNS_PRIME_BITS'd1098654767, `RNS_PRIME_BITS'd1477330056, `RNS_PRIME_BITS'd1569331694, `RNS_PRIME_BITS'd503094350 },
'{ `RNS_PRIME_BITS'd2014745094, `RNS_PRIME_BITS'd1203280856, `RNS_PRIME_BITS'd1874657457, `RNS_PRIME_BITS'd664236066, `RNS_PRIME_BITS'd1343163396, `RNS_PRIME_BITS'd349851856, `RNS_PRIME_BITS'd327986115, `RNS_PRIME_BITS'd1527009020, `RNS_PRIME_BITS'd1664893238, `RNS_PRIME_BITS'd2028124638 },
'{ `RNS_PRIME_BITS'd17214643, `RNS_PRIME_BITS'd1528026480, `RNS_PRIME_BITS'd707649348, `RNS_PRIME_BITS'd506168135, `RNS_PRIME_BITS'd623405378, `RNS_PRIME_BITS'd1082352090, `RNS_PRIME_BITS'd1990243254, `RNS_PRIME_BITS'd747636934, `RNS_PRIME_BITS'd1326828836, `RNS_PRIME_BITS'd1378524818 },
'{ `RNS_PRIME_BITS'd1873007184, `RNS_PRIME_BITS'd1982800586, `RNS_PRIME_BITS'd1616965474, `RNS_PRIME_BITS'd936503592, `RNS_PRIME_BITS'd265687623, `RNS_PRIME_BITS'd555195787, `RNS_PRIME_BITS'd703316243, `RNS_PRIME_BITS'd1230764655, `RNS_PRIME_BITS'd220437154, `RNS_PRIME_BITS'd1158294204 },
'{ `RNS_PRIME_BITS'd1171115647, `RNS_PRIME_BITS'd1636056387, `RNS_PRIME_BITS'd89367338, `RNS_PRIME_BITS'd1569217605, `RNS_PRIME_BITS'd148010597, `RNS_PRIME_BITS'd552135592, `RNS_PRIME_BITS'd1046145070, `RNS_PRIME_BITS'd1622489461, `RNS_PRIME_BITS'd627687042, `RNS_PRIME_BITS'd765167266 },
'{ `RNS_PRIME_BITS'd1810327907, `RNS_PRIME_BITS'd659636710, `RNS_PRIME_BITS'd527709368, `RNS_PRIME_BITS'd1981502868, `RNS_PRIME_BITS'd395782026, `RNS_PRIME_BITS'd1625981468, `RNS_PRIME_BITS'd263854684, `RNS_PRIME_BITS'd1651540472, `RNS_PRIME_BITS'd1368489211, `RNS_PRIME_BITS'd1257824607 }
};
parameter rns_residue_t y_q_TO_BBa[`B_BASIS_LEN +`Ba_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};


`define REG_NPOLY 12// how many polynomials can the register file store

// ---------------------------
// Operation/Control Types
// ---------------------------

// If you ever want to explicitly tag A vs B in code:
typedef enum logic [0:0] {
  POLY_A = 1'b0,
  POLY_B = 1'b1
} poly_sel_e;

typedef enum logic [1:0] {
    OP_CT_CT_ADD,
    OP_CT_PT_ADD,
    OP_CT_PT_MUL
} op_e;

typedef struct packed {
  op_e                          mode;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_b;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_b;
  logic [$clog2(`REG_NPOLY)-1:0]      out_a;
  logic [$clog2(`REG_NPOLY)-1:0]      out_b;
} operation;


`endif
