`ifndef TYPES_SVH
`define TYPES_SVH

// ---------------------------
// Basic data types
// ---------------------------

// NTT
`define BASE      32'd2
// Width of each RNS residue (one small prime)
`define RNS_PRIME_BITS 32
// RNS residues
typedef logic [`RNS_PRIME_BITS-1:0] rns_residue_t; 
typedef logic [(2*`RNS_PRIME_BITS)-1:0] wide_rns_residue_t;
// Vector / slot params
`define N_SLOTS   64
// moduli and RNS bases
`define t_MODULUS 257
`define q_BASIS_LEN 11
//`define q_MODULUS = 536101602793438606117677139878481445141305219292564418257989499598673136318603910408347407493377
parameter rns_residue_t q_BASIS [`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147492353, `RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193};
`define B_BASIS_LEN 10
//`define B_MODULUS = 2086194911538248702527219268311009200431885299167289996057309751033420854383242863211079351809
parameter rns_residue_t B_BASIS [`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147506433, `RNS_PRIME_BITS'd2147513089, `RNS_PRIME_BITS'd2147513857, `RNS_PRIME_BITS'd2147515649, `RNS_PRIME_BITS'd2147518721, `RNS_PRIME_BITS'd2147523841, `RNS_PRIME_BITS'd2147524097};
`define Ba_BASIS_LEN 10
//`define Ba_MODULUS = 2086476446457441129124572150314410036603537154987708995967124705067205076073473082954422397441
parameter rns_residue_t Ba_BASIS [`Ba_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147526401, `RNS_PRIME_BITS'd2147531777, `RNS_PRIME_BITS'd2147535617, `RNS_PRIME_BITS'd2147538433, `RNS_PRIME_BITS'd2147538689, `RNS_PRIME_BITS'd2147541761, `RNS_PRIME_BITS'd2147546113, `RNS_PRIME_BITS'd2147546881, `RNS_PRIME_BITS'd2147548673, `RNS_PRIME_BITS'd2147549953};
`define qBBa_BASIS_LEN 31
//`define qBBa_MODULUS = 2333541204753448940917127480778169670197024678706860035565116012612789108276505612899808761161753224723073709007431342423542638605605858321003804170268443281967101871649789313936832997411251353783868984682779840063476468468817175784888079498630244730925454530112323762437082863046913
parameter rns_residue_t qBBa_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147492353, `RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147506433, `RNS_PRIME_BITS'd2147513089, `RNS_PRIME_BITS'd2147513857, `RNS_PRIME_BITS'd2147515649, `RNS_PRIME_BITS'd2147518721, `RNS_PRIME_BITS'd2147523841, `RNS_PRIME_BITS'd2147524097, `RNS_PRIME_BITS'd2147526401, `RNS_PRIME_BITS'd2147531777, `RNS_PRIME_BITS'd2147535617, `RNS_PRIME_BITS'd2147538433, `RNS_PRIME_BITS'd2147538689, `RNS_PRIME_BITS'd2147541761, `RNS_PRIME_BITS'd2147546113, `RNS_PRIME_BITS'd2147546881, `RNS_PRIME_BITS'd2147548673, `RNS_PRIME_BITS'd2147549953};
// RNS integers
typedef rns_residue_t rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef rns_residue_t rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef rns_residue_t rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
/*typedef rns_residue_t rns_coef_qBBa_BASIS_t [`q_BASIS_LEN + `B_BASIS_LEN + `Ba_BASIS_LEN];*/
// Polynomials
typedef rns_int_q_BASIS_t q_BASIS_poly [`N_SLOTS];
typedef rns_int_B_BASIS_t B_BASIS_poly [`N_SLOTS];
typedef rns_int_Ba_BASIS_t Ba_BASIS_poly [`N_SLOTS];
/*typedef rns_coef_qBBA_BASIS_t qBBa_BASIS_poly [`N_SLOTS];*/
// wide RNS integers (each residue is double the length for mult)
typedef wide_rns_residue_t wide_rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
// wide Polynomials
typedef wide_rns_int_q_BASIS_t wide_q_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_B_BASIS_t wide_B_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_Ba_BASIS_t wide_Ba_BASIS_poly [`N_SLOTS];

// ---------------------------
// precalculated values
// ---------------------------
// Example constant “twist” factors (all 1s for now)
parameter rns_residue_t twist_factor   [`N_SLOTS] = '{default: '1};
parameter rns_residue_t untwist_factor [`N_SLOTS] = '{default: '1};

// fastBConv precalculated inverses
parameter rns_residue_t z_MOD_q [`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1065919626, `RNS_PRIME_BITS'd167960796, `RNS_PRIME_BITS'd20493556, `RNS_PRIME_BITS'd251993379, `RNS_PRIME_BITS'd574575462, `RNS_PRIME_BITS'd946908348, `RNS_PRIME_BITS'd907629872, `RNS_PRIME_BITS'd1497438013, `RNS_PRIME_BITS'd1737926542, `RNS_PRIME_BITS'd909409582};
parameter rns_residue_t z_MOD_B [`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd1692072777, `RNS_PRIME_BITS'd1095115435, `RNS_PRIME_BITS'd583606723, `RNS_PRIME_BITS'd2032025658, `RNS_PRIME_BITS'd394815268, `RNS_PRIME_BITS'd440518352, `RNS_PRIME_BITS'd1616527857, `RNS_PRIME_BITS'd1404316967, `RNS_PRIME_BITS'd961677545, `RNS_PRIME_BITS'd516873248};
parameter rns_residue_t y_q_TO_qBBa [`qBBa_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1181972137, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd25406470, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd225251055, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd708733459, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd626081157, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1145159656, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd2141619998, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd341559816, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd862367171, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd269122457 },
'{ `RNS_PRIME_BITS'd684423446, `RNS_PRIME_BITS'd204698767, `RNS_PRIME_BITS'd1405741688, `RNS_PRIME_BITS'd292426810, `RNS_PRIME_BITS'd649135386, `RNS_PRIME_BITS'd1045829233, `RNS_PRIME_BITS'd981025249, `RNS_PRIME_BITS'd494995369, `RNS_PRIME_BITS'd1816241534, `RNS_PRIME_BITS'd2046987670, `RNS_PRIME_BITS'd1979981476 },
'{ `RNS_PRIME_BITS'd906641143, `RNS_PRIME_BITS'd1415238335, `RNS_PRIME_BITS'd1263671982, `RNS_PRIME_BITS'd1171151273, `RNS_PRIME_BITS'd194982496, `RNS_PRIME_BITS'd885154054, `RNS_PRIME_BITS'd520252441, `RNS_PRIME_BITS'd2102695851, `RNS_PRIME_BITS'd1854128422, `RNS_PRIME_BITS'd1365954298, `RNS_PRIME_BITS'd584947488 },
'{ `RNS_PRIME_BITS'd1468203946, `RNS_PRIME_BITS'd1481404946, `RNS_PRIME_BITS'd1609922880, `RNS_PRIME_BITS'd1341334258, `RNS_PRIME_BITS'd1330494182, `RNS_PRIME_BITS'd824735172, `RNS_PRIME_BITS'd394332974, `RNS_PRIME_BITS'd1560369477, `RNS_PRIME_BITS'd738867587, `RNS_PRIME_BITS'd1237102758, `RNS_PRIME_BITS'd266443486 },
'{ `RNS_PRIME_BITS'd1418389148, `RNS_PRIME_BITS'd270198595, `RNS_PRIME_BITS'd1276905103, `RNS_PRIME_BITS'd1847640359, `RNS_PRIME_BITS'd453784804, `RNS_PRIME_BITS'd1403544338, `RNS_PRIME_BITS'd1747685001, `RNS_PRIME_BITS'd1575406910, `RNS_PRIME_BITS'd1238219428, `RNS_PRIME_BITS'd406303773, `RNS_PRIME_BITS'd319243640 },
'{ `RNS_PRIME_BITS'd98660650, `RNS_PRIME_BITS'd382332231, `RNS_PRIME_BITS'd1232241863, `RNS_PRIME_BITS'd1339301824, `RNS_PRIME_BITS'd773056655, `RNS_PRIME_BITS'd533377063, `RNS_PRIME_BITS'd352136881, `RNS_PRIME_BITS'd1950455605, `RNS_PRIME_BITS'd608500593, `RNS_PRIME_BITS'd1298548779, `RNS_PRIME_BITS'd1337898742 },
'{ `RNS_PRIME_BITS'd1792684747, `RNS_PRIME_BITS'd573070289, `RNS_PRIME_BITS'd1500502820, `RNS_PRIME_BITS'd1933930544, `RNS_PRIME_BITS'd202429986, `RNS_PRIME_BITS'd1609483297, `RNS_PRIME_BITS'd205823311, `RNS_PRIME_BITS'd1072516210, `RNS_PRIME_BITS'd2001103785, `RNS_PRIME_BITS'd1329490615, `RNS_PRIME_BITS'd1119039461 },
'{ `RNS_PRIME_BITS'd951706160, `RNS_PRIME_BITS'd292317085, `RNS_PRIME_BITS'd31185556, `RNS_PRIME_BITS'd1704940567, `RNS_PRIME_BITS'd920960039, `RNS_PRIME_BITS'd1433469121, `RNS_PRIME_BITS'd757419291, `RNS_PRIME_BITS'd675648917, `RNS_PRIME_BITS'd841576990, `RNS_PRIME_BITS'd2030299916, `RNS_PRIME_BITS'd162267491 },
'{ `RNS_PRIME_BITS'd1832276929, `RNS_PRIME_BITS'd1668659698, `RNS_PRIME_BITS'd1999427244, `RNS_PRIME_BITS'd1340362480, `RNS_PRIME_BITS'd1749989777, `RNS_PRIME_BITS'd498252843, `RNS_PRIME_BITS'd1324247774, `RNS_PRIME_BITS'd573351343, `RNS_PRIME_BITS'd2006599164, `RNS_PRIME_BITS'd355470826, `RNS_PRIME_BITS'd851622145 },
'{ `RNS_PRIME_BITS'd1368158453, `RNS_PRIME_BITS'd1057377784, `RNS_PRIME_BITS'd1982467647, `RNS_PRIME_BITS'd1477457381, `RNS_PRIME_BITS'd389718782, `RNS_PRIME_BITS'd1035655701, `RNS_PRIME_BITS'd146409306, `RNS_PRIME_BITS'd1419154533, `RNS_PRIME_BITS'd2001519893, `RNS_PRIME_BITS'd1685170863, `RNS_PRIME_BITS'd2074298371 },
'{ `RNS_PRIME_BITS'd322502136, `RNS_PRIME_BITS'd1511774222, `RNS_PRIME_BITS'd615033910, `RNS_PRIME_BITS'd1032913238, `RNS_PRIME_BITS'd1412879797, `RNS_PRIME_BITS'd1416984709, `RNS_PRIME_BITS'd1917372184, `RNS_PRIME_BITS'd1707427060, `RNS_PRIME_BITS'd1616633336, `RNS_PRIME_BITS'd1312078978, `RNS_PRIME_BITS'd2143938115 },
'{ `RNS_PRIME_BITS'd1739800961, `RNS_PRIME_BITS'd1466703262, `RNS_PRIME_BITS'd698484285, `RNS_PRIME_BITS'd1183868308, `RNS_PRIME_BITS'd1591117221, `RNS_PRIME_BITS'd1674272937, `RNS_PRIME_BITS'd759615877, `RNS_PRIME_BITS'd1009347551, `RNS_PRIME_BITS'd553304063, `RNS_PRIME_BITS'd1479835385, `RNS_PRIME_BITS'd1395721083 },
'{ `RNS_PRIME_BITS'd1778336261, `RNS_PRIME_BITS'd648741787, `RNS_PRIME_BITS'd941020410, `RNS_PRIME_BITS'd1007056930, `RNS_PRIME_BITS'd1043677182, `RNS_PRIME_BITS'd1425015806, `RNS_PRIME_BITS'd367581824, `RNS_PRIME_BITS'd554124327, `RNS_PRIME_BITS'd390555688, `RNS_PRIME_BITS'd1815322513, `RNS_PRIME_BITS'd1594244359 },
'{ `RNS_PRIME_BITS'd756715838, `RNS_PRIME_BITS'd479599688, `RNS_PRIME_BITS'd1528095740, `RNS_PRIME_BITS'd1349581192, `RNS_PRIME_BITS'd1680905314, `RNS_PRIME_BITS'd1116825851, `RNS_PRIME_BITS'd880597572, `RNS_PRIME_BITS'd960310028, `RNS_PRIME_BITS'd2064989836, `RNS_PRIME_BITS'd2104701179, `RNS_PRIME_BITS'd1351112918 },
'{ `RNS_PRIME_BITS'd1760592201, `RNS_PRIME_BITS'd1898972358, `RNS_PRIME_BITS'd1309712124, `RNS_PRIME_BITS'd1433096384, `RNS_PRIME_BITS'd387480417, `RNS_PRIME_BITS'd2093398215, `RNS_PRIME_BITS'd1841149906, `RNS_PRIME_BITS'd314258125, `RNS_PRIME_BITS'd447978224, `RNS_PRIME_BITS'd970406200, `RNS_PRIME_BITS'd2088476377 },
'{ `RNS_PRIME_BITS'd874133271, `RNS_PRIME_BITS'd97609305, `RNS_PRIME_BITS'd2093146792, `RNS_PRIME_BITS'd788311714, `RNS_PRIME_BITS'd678725287, `RNS_PRIME_BITS'd886081750, `RNS_PRIME_BITS'd1726158361, `RNS_PRIME_BITS'd1223252937, `RNS_PRIME_BITS'd1703980449, `RNS_PRIME_BITS'd468894801, `RNS_PRIME_BITS'd8812854 },
'{ `RNS_PRIME_BITS'd513828569, `RNS_PRIME_BITS'd1733376001, `RNS_PRIME_BITS'd276737436, `RNS_PRIME_BITS'd783417692, `RNS_PRIME_BITS'd427481431, `RNS_PRIME_BITS'd2087538087, `RNS_PRIME_BITS'd1662191261, `RNS_PRIME_BITS'd1247267656, `RNS_PRIME_BITS'd1567910359, `RNS_PRIME_BITS'd1629834561, `RNS_PRIME_BITS'd1720536357 },
'{ `RNS_PRIME_BITS'd1116386599, `RNS_PRIME_BITS'd511421869, `RNS_PRIME_BITS'd131462801, `RNS_PRIME_BITS'd81649043, `RNS_PRIME_BITS'd1454019614, `RNS_PRIME_BITS'd16673857, `RNS_PRIME_BITS'd818230176, `RNS_PRIME_BITS'd1217263563, `RNS_PRIME_BITS'd1198657912, `RNS_PRIME_BITS'd1009787849, `RNS_PRIME_BITS'd1504719155 },
'{ `RNS_PRIME_BITS'd2039477880, `RNS_PRIME_BITS'd1398231506, `RNS_PRIME_BITS'd1983511237, `RNS_PRIME_BITS'd368961275, `RNS_PRIME_BITS'd52877229, `RNS_PRIME_BITS'd1144504988, `RNS_PRIME_BITS'd339508547, `RNS_PRIME_BITS'd2080271213, `RNS_PRIME_BITS'd1983734146, `RNS_PRIME_BITS'd2034965627, `RNS_PRIME_BITS'd515360951 },
'{ `RNS_PRIME_BITS'd472567105, `RNS_PRIME_BITS'd1909213356, `RNS_PRIME_BITS'd1440608399, `RNS_PRIME_BITS'd1486366436, `RNS_PRIME_BITS'd1887546509, `RNS_PRIME_BITS'd586017197, `RNS_PRIME_BITS'd1961555240, `RNS_PRIME_BITS'd1084140746, `RNS_PRIME_BITS'd1432036558, `RNS_PRIME_BITS'd1950773012, `RNS_PRIME_BITS'd1414585043 },
'{ `RNS_PRIME_BITS'd755457487, `RNS_PRIME_BITS'd1733544464, `RNS_PRIME_BITS'd215223763, `RNS_PRIME_BITS'd776094764, `RNS_PRIME_BITS'd1341813263, `RNS_PRIME_BITS'd395678378, `RNS_PRIME_BITS'd608364884, `RNS_PRIME_BITS'd377100389, `RNS_PRIME_BITS'd264252957, `RNS_PRIME_BITS'd1655795893, `RNS_PRIME_BITS'd1651112521 }
};
parameter rns_residue_t y_B_TO_Ba[`Ba_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd536926448, `RNS_PRIME_BITS'd997114948, `RNS_PRIME_BITS'd2119023736, `RNS_PRIME_BITS'd20715414, `RNS_PRIME_BITS'd31073121, `RNS_PRIME_BITS'd1216306431, `RNS_PRIME_BITS'd345260969, `RNS_PRIME_BITS'd1342375917, `RNS_PRIME_BITS'd1879601350, `RNS_PRIME_BITS'd179533588 },
'{ `RNS_PRIME_BITS'd736010931, `RNS_PRIME_BITS'd692161079, `RNS_PRIME_BITS'd814390359, `RNS_PRIME_BITS'd1466622767, `RNS_PRIME_BITS'd1665380882, `RNS_PRIME_BITS'd2104902653, `RNS_PRIME_BITS'd1384322158, `RNS_PRIME_BITS'd1962695816, `RNS_PRIME_BITS'd1289245060, `RNS_PRIME_BITS'd2048063821 },
'{ `RNS_PRIME_BITS'd1606987083, `RNS_PRIME_BITS'd350190383, `RNS_PRIME_BITS'd1222316619, `RNS_PRIME_BITS'd263587925, `RNS_PRIME_BITS'd1854502633, `RNS_PRIME_BITS'd606169172, `RNS_PRIME_BITS'd2037194365, `RNS_PRIME_BITS'd1040979766, `RNS_PRIME_BITS'd746610754, `RNS_PRIME_BITS'd2099446488 },
'{ `RNS_PRIME_BITS'd728466737, `RNS_PRIME_BITS'd635106757, `RNS_PRIME_BITS'd334346405, `RNS_PRIME_BITS'd1493862730, `RNS_PRIME_BITS'd1582498012, `RNS_PRIME_BITS'd1900393379, `RNS_PRIME_BITS'd119490896, `RNS_PRIME_BITS'd1114266687, `RNS_PRIME_BITS'd261925730, `RNS_PRIME_BITS'd189905174 },
'{ `RNS_PRIME_BITS'd2060710709, `RNS_PRIME_BITS'd1002320634, `RNS_PRIME_BITS'd958977095, `RNS_PRIME_BITS'd1217103627, `RNS_PRIME_BITS'd1146993606, `RNS_PRIME_BITS'd1758096562, `RNS_PRIME_BITS'd1274437340, `RNS_PRIME_BITS'd809723488, `RNS_PRIME_BITS'd2051628241, `RNS_PRIME_BITS'd1560156076 },
'{ `RNS_PRIME_BITS'd635786634, `RNS_PRIME_BITS'd1455243434, `RNS_PRIME_BITS'd332022673, `RNS_PRIME_BITS'd59280119, `RNS_PRIME_BITS'd1798744776, `RNS_PRIME_BITS'd1749740423, `RNS_PRIME_BITS'd2101418289, `RNS_PRIME_BITS'd1952099042, `RNS_PRIME_BITS'd1589466585, `RNS_PRIME_BITS'd118560238 },
'{ `RNS_PRIME_BITS'd1069408896, `RNS_PRIME_BITS'd490983615, `RNS_PRIME_BITS'd1765883527, `RNS_PRIME_BITS'd1546369328, `RNS_PRIME_BITS'd1891335954, `RNS_PRIME_BITS'd709198555, `RNS_PRIME_BITS'd877242359, `RNS_PRIME_BITS'd1136188875, `RNS_PRIME_BITS'd2063861548, `RNS_PRIME_BITS'd689457818 },
'{ `RNS_PRIME_BITS'd472953696, `RNS_PRIME_BITS'd1020895029, `RNS_PRIME_BITS'd1196514381, `RNS_PRIME_BITS'd1344864532, `RNS_PRIME_BITS'd893913131, `RNS_PRIME_BITS'd1713789020, `RNS_PRIME_BITS'd1389652938, `RNS_PRIME_BITS'd643186381, `RNS_PRIME_BITS'd1024733008, `RNS_PRIME_BITS'd215835694 },
'{ `RNS_PRIME_BITS'd516845021, `RNS_PRIME_BITS'd163468955, `RNS_PRIME_BITS'd1181920865, `RNS_PRIME_BITS'd775913513, `RNS_PRIME_BITS'd1817147861, `RNS_PRIME_BITS'd1620370019, `RNS_PRIME_BITS'd1292105471, `RNS_PRIME_BITS'd1699955862, `RNS_PRIME_BITS'd279288062, `RNS_PRIME_BITS'd326937910 },
'{ `RNS_PRIME_BITS'd609874074, `RNS_PRIME_BITS'd1436624771, `RNS_PRIME_BITS'd2064246923, `RNS_PRIME_BITS'd1930080170, `RNS_PRIME_BITS'd71362749, `RNS_PRIME_BITS'd941039597, `RNS_PRIME_BITS'd653642046, `RNS_PRIME_BITS'd858757654, `RNS_PRIME_BITS'd353400346, `RNS_PRIME_BITS'd37956297 }
};
parameter rns_residue_t y_B_TO_q[`q_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd73 },
'{ `RNS_PRIME_BITS'd70868141, `RNS_PRIME_BITS'd416970811, `RNS_PRIME_BITS'd987541071, `RNS_PRIME_BITS'd1472384924, `RNS_PRIME_BITS'd544473269, `RNS_PRIME_BITS'd1104288693, `RNS_PRIME_BITS'd360533383, `RNS_PRIME_BITS'd1855585819, `RNS_PRIME_BITS'd854144882, `RNS_PRIME_BITS'd1316711014 },
'{ `RNS_PRIME_BITS'd629451863, `RNS_PRIME_BITS'd1573926589, `RNS_PRIME_BITS'd782449585, `RNS_PRIME_BITS'd837933943, `RNS_PRIME_BITS'd1069373815, `RNS_PRIME_BITS'd679901823, `RNS_PRIME_BITS'd801302253, `RNS_PRIME_BITS'd533230691, `RNS_PRIME_BITS'd858658087, `RNS_PRIME_BITS'd2018021427 },
'{ `RNS_PRIME_BITS'd1358250437, `RNS_PRIME_BITS'd101977895, `RNS_PRIME_BITS'd580470523, `RNS_PRIME_BITS'd1405916185, `RNS_PRIME_BITS'd945265442, `RNS_PRIME_BITS'd1959038865, `RNS_PRIME_BITS'd221448123, `RNS_PRIME_BITS'd843549711, `RNS_PRIME_BITS'd1950178610, `RNS_PRIME_BITS'd1677430563 },
'{ `RNS_PRIME_BITS'd1619523558, `RNS_PRIME_BITS'd378303593, `RNS_PRIME_BITS'd1540620734, `RNS_PRIME_BITS'd321156193, `RNS_PRIME_BITS'd1397508539, `RNS_PRIME_BITS'd923878783, `RNS_PRIME_BITS'd1092067346, `RNS_PRIME_BITS'd411984063, `RNS_PRIME_BITS'd2081306367, `RNS_PRIME_BITS'd1206893468 },
'{ `RNS_PRIME_BITS'd1932818330, `RNS_PRIME_BITS'd1856095313, `RNS_PRIME_BITS'd726878279, `RNS_PRIME_BITS'd1999144769, `RNS_PRIME_BITS'd190904923, `RNS_PRIME_BITS'd1334529222, `RNS_PRIME_BITS'd1231873128, `RNS_PRIME_BITS'd2089127064, `RNS_PRIME_BITS'd492362912, `RNS_PRIME_BITS'd142022509 },
'{ `RNS_PRIME_BITS'd1582143434, `RNS_PRIME_BITS'd359870278, `RNS_PRIME_BITS'd142671376, `RNS_PRIME_BITS'd179935139, `RNS_PRIME_BITS'd1356264469, `RNS_PRIME_BITS'd479293904, `RNS_PRIME_BITS'd966958127, `RNS_PRIME_BITS'd979521442, `RNS_PRIME_BITS'd396486594, `RNS_PRIME_BITS'd1440820496 },
'{ `RNS_PRIME_BITS'd1767412547, `RNS_PRIME_BITS'd1549723359, `RNS_PRIME_BITS'd1033148906, `RNS_PRIME_BITS'd345182914, `RNS_PRIME_BITS'd969984052, `RNS_PRIME_BITS'd106717785, `RNS_PRIME_BITS'd1234837791, `RNS_PRIME_BITS'd1259187251, `RNS_PRIME_BITS'd71145190, `RNS_PRIME_BITS'd1526470325 },
'{ `RNS_PRIME_BITS'd772904767, `RNS_PRIME_BITS'd2013787051, `RNS_PRIME_BITS'd1323988339, `RNS_PRIME_BITS'd1235013803, `RNS_PRIME_BITS'd480291155, `RNS_PRIME_BITS'd2114971379, `RNS_PRIME_BITS'd1640560963, `RNS_PRIME_BITS'd1359601648, `RNS_PRIME_BITS'd814894112, `RNS_PRIME_BITS'd1448226857 },
'{ `RNS_PRIME_BITS'd572041956, `RNS_PRIME_BITS'd190680652, `RNS_PRIME_BITS'd2092311774, `RNS_PRIME_BITS'd1295240622, `RNS_PRIME_BITS'd926324836, `RNS_PRIME_BITS'd191516735, `RNS_PRIME_BITS'd697437258, `RNS_PRIME_BITS'd1463443896, `RNS_PRIME_BITS'd1978270708, `RNS_PRIME_BITS'd1766980370 },
'{ `RNS_PRIME_BITS'd812796495, `RNS_PRIME_BITS'd1178720511, `RNS_PRIME_BITS'd370036586, `RNS_PRIME_BITS'd1940018906, `RNS_PRIME_BITS'd1501147245, `RNS_PRIME_BITS'd969032975, `RNS_PRIME_BITS'd455932005, `RNS_PRIME_BITS'd1662734482, `RNS_PRIME_BITS'd1275283793, `RNS_PRIME_BITS'd554319144 }
};
parameter rns_residue_t y_q_TO_BBa[`B_BASIS_LEN +`Ba_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd684423446, `RNS_PRIME_BITS'd204698767, `RNS_PRIME_BITS'd1405741688, `RNS_PRIME_BITS'd292426810, `RNS_PRIME_BITS'd649135386, `RNS_PRIME_BITS'd1045829233, `RNS_PRIME_BITS'd981025249, `RNS_PRIME_BITS'd494995369, `RNS_PRIME_BITS'd1816241534, `RNS_PRIME_BITS'd2046987670, `RNS_PRIME_BITS'd1979981476 },
'{ `RNS_PRIME_BITS'd906641143, `RNS_PRIME_BITS'd1415238335, `RNS_PRIME_BITS'd1263671982, `RNS_PRIME_BITS'd1171151273, `RNS_PRIME_BITS'd194982496, `RNS_PRIME_BITS'd885154054, `RNS_PRIME_BITS'd520252441, `RNS_PRIME_BITS'd2102695851, `RNS_PRIME_BITS'd1854128422, `RNS_PRIME_BITS'd1365954298, `RNS_PRIME_BITS'd584947488 },
'{ `RNS_PRIME_BITS'd1468203946, `RNS_PRIME_BITS'd1481404946, `RNS_PRIME_BITS'd1609922880, `RNS_PRIME_BITS'd1341334258, `RNS_PRIME_BITS'd1330494182, `RNS_PRIME_BITS'd824735172, `RNS_PRIME_BITS'd394332974, `RNS_PRIME_BITS'd1560369477, `RNS_PRIME_BITS'd738867587, `RNS_PRIME_BITS'd1237102758, `RNS_PRIME_BITS'd266443486 },
'{ `RNS_PRIME_BITS'd1418389148, `RNS_PRIME_BITS'd270198595, `RNS_PRIME_BITS'd1276905103, `RNS_PRIME_BITS'd1847640359, `RNS_PRIME_BITS'd453784804, `RNS_PRIME_BITS'd1403544338, `RNS_PRIME_BITS'd1747685001, `RNS_PRIME_BITS'd1575406910, `RNS_PRIME_BITS'd1238219428, `RNS_PRIME_BITS'd406303773, `RNS_PRIME_BITS'd319243640 },
'{ `RNS_PRIME_BITS'd98660650, `RNS_PRIME_BITS'd382332231, `RNS_PRIME_BITS'd1232241863, `RNS_PRIME_BITS'd1339301824, `RNS_PRIME_BITS'd773056655, `RNS_PRIME_BITS'd533377063, `RNS_PRIME_BITS'd352136881, `RNS_PRIME_BITS'd1950455605, `RNS_PRIME_BITS'd608500593, `RNS_PRIME_BITS'd1298548779, `RNS_PRIME_BITS'd1337898742 },
'{ `RNS_PRIME_BITS'd1792684747, `RNS_PRIME_BITS'd573070289, `RNS_PRIME_BITS'd1500502820, `RNS_PRIME_BITS'd1933930544, `RNS_PRIME_BITS'd202429986, `RNS_PRIME_BITS'd1609483297, `RNS_PRIME_BITS'd205823311, `RNS_PRIME_BITS'd1072516210, `RNS_PRIME_BITS'd2001103785, `RNS_PRIME_BITS'd1329490615, `RNS_PRIME_BITS'd1119039461 },
'{ `RNS_PRIME_BITS'd951706160, `RNS_PRIME_BITS'd292317085, `RNS_PRIME_BITS'd31185556, `RNS_PRIME_BITS'd1704940567, `RNS_PRIME_BITS'd920960039, `RNS_PRIME_BITS'd1433469121, `RNS_PRIME_BITS'd757419291, `RNS_PRIME_BITS'd675648917, `RNS_PRIME_BITS'd841576990, `RNS_PRIME_BITS'd2030299916, `RNS_PRIME_BITS'd162267491 },
'{ `RNS_PRIME_BITS'd1832276929, `RNS_PRIME_BITS'd1668659698, `RNS_PRIME_BITS'd1999427244, `RNS_PRIME_BITS'd1340362480, `RNS_PRIME_BITS'd1749989777, `RNS_PRIME_BITS'd498252843, `RNS_PRIME_BITS'd1324247774, `RNS_PRIME_BITS'd573351343, `RNS_PRIME_BITS'd2006599164, `RNS_PRIME_BITS'd355470826, `RNS_PRIME_BITS'd851622145 },
'{ `RNS_PRIME_BITS'd1368158453, `RNS_PRIME_BITS'd1057377784, `RNS_PRIME_BITS'd1982467647, `RNS_PRIME_BITS'd1477457381, `RNS_PRIME_BITS'd389718782, `RNS_PRIME_BITS'd1035655701, `RNS_PRIME_BITS'd146409306, `RNS_PRIME_BITS'd1419154533, `RNS_PRIME_BITS'd2001519893, `RNS_PRIME_BITS'd1685170863, `RNS_PRIME_BITS'd2074298371 },
'{ `RNS_PRIME_BITS'd322502136, `RNS_PRIME_BITS'd1511774222, `RNS_PRIME_BITS'd615033910, `RNS_PRIME_BITS'd1032913238, `RNS_PRIME_BITS'd1412879797, `RNS_PRIME_BITS'd1416984709, `RNS_PRIME_BITS'd1917372184, `RNS_PRIME_BITS'd1707427060, `RNS_PRIME_BITS'd1616633336, `RNS_PRIME_BITS'd1312078978, `RNS_PRIME_BITS'd2143938115 },
'{ `RNS_PRIME_BITS'd1739800961, `RNS_PRIME_BITS'd1466703262, `RNS_PRIME_BITS'd698484285, `RNS_PRIME_BITS'd1183868308, `RNS_PRIME_BITS'd1591117221, `RNS_PRIME_BITS'd1674272937, `RNS_PRIME_BITS'd759615877, `RNS_PRIME_BITS'd1009347551, `RNS_PRIME_BITS'd553304063, `RNS_PRIME_BITS'd1479835385, `RNS_PRIME_BITS'd1395721083 },
'{ `RNS_PRIME_BITS'd1778336261, `RNS_PRIME_BITS'd648741787, `RNS_PRIME_BITS'd941020410, `RNS_PRIME_BITS'd1007056930, `RNS_PRIME_BITS'd1043677182, `RNS_PRIME_BITS'd1425015806, `RNS_PRIME_BITS'd367581824, `RNS_PRIME_BITS'd554124327, `RNS_PRIME_BITS'd390555688, `RNS_PRIME_BITS'd1815322513, `RNS_PRIME_BITS'd1594244359 },
'{ `RNS_PRIME_BITS'd756715838, `RNS_PRIME_BITS'd479599688, `RNS_PRIME_BITS'd1528095740, `RNS_PRIME_BITS'd1349581192, `RNS_PRIME_BITS'd1680905314, `RNS_PRIME_BITS'd1116825851, `RNS_PRIME_BITS'd880597572, `RNS_PRIME_BITS'd960310028, `RNS_PRIME_BITS'd2064989836, `RNS_PRIME_BITS'd2104701179, `RNS_PRIME_BITS'd1351112918 },
'{ `RNS_PRIME_BITS'd1760592201, `RNS_PRIME_BITS'd1898972358, `RNS_PRIME_BITS'd1309712124, `RNS_PRIME_BITS'd1433096384, `RNS_PRIME_BITS'd387480417, `RNS_PRIME_BITS'd2093398215, `RNS_PRIME_BITS'd1841149906, `RNS_PRIME_BITS'd314258125, `RNS_PRIME_BITS'd447978224, `RNS_PRIME_BITS'd970406200, `RNS_PRIME_BITS'd2088476377 },
'{ `RNS_PRIME_BITS'd874133271, `RNS_PRIME_BITS'd97609305, `RNS_PRIME_BITS'd2093146792, `RNS_PRIME_BITS'd788311714, `RNS_PRIME_BITS'd678725287, `RNS_PRIME_BITS'd886081750, `RNS_PRIME_BITS'd1726158361, `RNS_PRIME_BITS'd1223252937, `RNS_PRIME_BITS'd1703980449, `RNS_PRIME_BITS'd468894801, `RNS_PRIME_BITS'd8812854 },
'{ `RNS_PRIME_BITS'd513828569, `RNS_PRIME_BITS'd1733376001, `RNS_PRIME_BITS'd276737436, `RNS_PRIME_BITS'd783417692, `RNS_PRIME_BITS'd427481431, `RNS_PRIME_BITS'd2087538087, `RNS_PRIME_BITS'd1662191261, `RNS_PRIME_BITS'd1247267656, `RNS_PRIME_BITS'd1567910359, `RNS_PRIME_BITS'd1629834561, `RNS_PRIME_BITS'd1720536357 },
'{ `RNS_PRIME_BITS'd1116386599, `RNS_PRIME_BITS'd511421869, `RNS_PRIME_BITS'd131462801, `RNS_PRIME_BITS'd81649043, `RNS_PRIME_BITS'd1454019614, `RNS_PRIME_BITS'd16673857, `RNS_PRIME_BITS'd818230176, `RNS_PRIME_BITS'd1217263563, `RNS_PRIME_BITS'd1198657912, `RNS_PRIME_BITS'd1009787849, `RNS_PRIME_BITS'd1504719155 },
'{ `RNS_PRIME_BITS'd2039477880, `RNS_PRIME_BITS'd1398231506, `RNS_PRIME_BITS'd1983511237, `RNS_PRIME_BITS'd368961275, `RNS_PRIME_BITS'd52877229, `RNS_PRIME_BITS'd1144504988, `RNS_PRIME_BITS'd339508547, `RNS_PRIME_BITS'd2080271213, `RNS_PRIME_BITS'd1983734146, `RNS_PRIME_BITS'd2034965627, `RNS_PRIME_BITS'd515360951 },
'{ `RNS_PRIME_BITS'd472567105, `RNS_PRIME_BITS'd1909213356, `RNS_PRIME_BITS'd1440608399, `RNS_PRIME_BITS'd1486366436, `RNS_PRIME_BITS'd1887546509, `RNS_PRIME_BITS'd586017197, `RNS_PRIME_BITS'd1961555240, `RNS_PRIME_BITS'd1084140746, `RNS_PRIME_BITS'd1432036558, `RNS_PRIME_BITS'd1950773012, `RNS_PRIME_BITS'd1414585043 },
'{ `RNS_PRIME_BITS'd755457487, `RNS_PRIME_BITS'd1733544464, `RNS_PRIME_BITS'd215223763, `RNS_PRIME_BITS'd776094764, `RNS_PRIME_BITS'd1341813263, `RNS_PRIME_BITS'd395678378, `RNS_PRIME_BITS'd608364884, `RNS_PRIME_BITS'd377100389, `RNS_PRIME_BITS'd264252957, `RNS_PRIME_BITS'd1655795893, `RNS_PRIME_BITS'd1651112521 }
};


`define REG_NPOLY 12// how many polynomials can the register file store

// ---------------------------
// Operation/Control Types
// ---------------------------

// If you ever want to explicitly tag A vs B in code:
typedef enum logic [0:0] {
  POLY_A = 1'b0,
  POLY_B = 1'b1
} poly_sel_e;

typedef enum logic [1:0] {
    OP_CT_CT_ADD,
    OP_CT_PT_ADD,
    OP_CT_PT_MUL
} op_e;

typedef struct packed {
  op_e                          mode;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_b;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_b;
  logic [$clog2(`REG_NPOLY)-1:0]      out_a;
  logic [$clog2(`REG_NPOLY)-1:0]      out_b;
} operation;


`endif
