`include "types.svh"

`ifndef CTEXAMPLES_SVH
`define CTEXAMPLES_SVH

const rns_residue_t A1__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1007849158, `RNS_PRIME_BITS'd344623035, `RNS_PRIME_BITS'd974553355, `RNS_PRIME_BITS'd252232956, `RNS_PRIME_BITS'd1591552870, `RNS_PRIME_BITS'd1997619035, `RNS_PRIME_BITS'd168382023, `RNS_PRIME_BITS'd978517921, `RNS_PRIME_BITS'd225318580, `RNS_PRIME_BITS'd108420664},
    '{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd1228814435, `RNS_PRIME_BITS'd151413131, `RNS_PRIME_BITS'd2050222428, `RNS_PRIME_BITS'd1413564231, `RNS_PRIME_BITS'd439481772, `RNS_PRIME_BITS'd444027837, `RNS_PRIME_BITS'd985258507, `RNS_PRIME_BITS'd583611165, `RNS_PRIME_BITS'd2035531980, `RNS_PRIME_BITS'd386692334},
    '{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd128486397, `RNS_PRIME_BITS'd1816285854, `RNS_PRIME_BITS'd863587800, `RNS_PRIME_BITS'd267914966, `RNS_PRIME_BITS'd1697223387, `RNS_PRIME_BITS'd1705853764, `RNS_PRIME_BITS'd775183607, `RNS_PRIME_BITS'd1128390963, `RNS_PRIME_BITS'd380101658, `RNS_PRIME_BITS'd1930921843},
    '{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd135710087, `RNS_PRIME_BITS'd1425278094, `RNS_PRIME_BITS'd1559673485, `RNS_PRIME_BITS'd176413468, `RNS_PRIME_BITS'd136727317, `RNS_PRIME_BITS'd1385941432, `RNS_PRIME_BITS'd1576270542, `RNS_PRIME_BITS'd71341352, `RNS_PRIME_BITS'd2081847665, `RNS_PRIME_BITS'd475256072},
    '{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd717104875, `RNS_PRIME_BITS'd2051774700, `RNS_PRIME_BITS'd368829184, `RNS_PRIME_BITS'd6013804, `RNS_PRIME_BITS'd383335523, `RNS_PRIME_BITS'd965384056, `RNS_PRIME_BITS'd1828281782, `RNS_PRIME_BITS'd407992677, `RNS_PRIME_BITS'd839636323, `RNS_PRIME_BITS'd1460582641},
    '{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd238512322, `RNS_PRIME_BITS'd2095782834, `RNS_PRIME_BITS'd1926466631, `RNS_PRIME_BITS'd348242689, `RNS_PRIME_BITS'd1452579508, `RNS_PRIME_BITS'd2076181866, `RNS_PRIME_BITS'd946667019, `RNS_PRIME_BITS'd248454984, `RNS_PRIME_BITS'd2108208234, `RNS_PRIME_BITS'd1417627426},
    '{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd2072819984, `RNS_PRIME_BITS'd1872956090, `RNS_PRIME_BITS'd534439250, `RNS_PRIME_BITS'd461321156, `RNS_PRIME_BITS'd1648784831, `RNS_PRIME_BITS'd1125878975, `RNS_PRIME_BITS'd562094147, `RNS_PRIME_BITS'd1584847967, `RNS_PRIME_BITS'd2030964712, `RNS_PRIME_BITS'd362752790},
    '{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1457932833, `RNS_PRIME_BITS'd1554698931, `RNS_PRIME_BITS'd136975177, `RNS_PRIME_BITS'd1209489831, `RNS_PRIME_BITS'd1234868194, `RNS_PRIME_BITS'd1474258431, `RNS_PRIME_BITS'd1725337056, `RNS_PRIME_BITS'd1411870778, `RNS_PRIME_BITS'd2058986111, `RNS_PRIME_BITS'd157537645},
    '{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd771191296, `RNS_PRIME_BITS'd1929166853, `RNS_PRIME_BITS'd220566812, `RNS_PRIME_BITS'd1515595715, `RNS_PRIME_BITS'd1047050759, `RNS_PRIME_BITS'd262115771, `RNS_PRIME_BITS'd1924947401, `RNS_PRIME_BITS'd512489747, `RNS_PRIME_BITS'd580532616, `RNS_PRIME_BITS'd1945613104},
    '{`RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd1929758221, `RNS_PRIME_BITS'd1996127246, `RNS_PRIME_BITS'd937804862, `RNS_PRIME_BITS'd1288253295, `RNS_PRIME_BITS'd1076311145, `RNS_PRIME_BITS'd144918156, `RNS_PRIME_BITS'd1842504095, `RNS_PRIME_BITS'd1278919215, `RNS_PRIME_BITS'd556241807, `RNS_PRIME_BITS'd100699118},
    '{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1661095827, `RNS_PRIME_BITS'd20449632, `RNS_PRIME_BITS'd1121730000, `RNS_PRIME_BITS'd361938300, `RNS_PRIME_BITS'd1772251391, `RNS_PRIME_BITS'd254315466, `RNS_PRIME_BITS'd438135027, `RNS_PRIME_BITS'd876666992, `RNS_PRIME_BITS'd798295796, `RNS_PRIME_BITS'd1458298158},
    '{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd916253055, `RNS_PRIME_BITS'd108274752, `RNS_PRIME_BITS'd1697816182, `RNS_PRIME_BITS'd903388280, `RNS_PRIME_BITS'd1716351348, `RNS_PRIME_BITS'd547309949, `RNS_PRIME_BITS'd1021283545, `RNS_PRIME_BITS'd1558943094, `RNS_PRIME_BITS'd38353636, `RNS_PRIME_BITS'd292512990},
    '{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1132664726, `RNS_PRIME_BITS'd1787992750, `RNS_PRIME_BITS'd1099387607, `RNS_PRIME_BITS'd1306070432, `RNS_PRIME_BITS'd1905096779, `RNS_PRIME_BITS'd1508222052, `RNS_PRIME_BITS'd325083905, `RNS_PRIME_BITS'd3522864, `RNS_PRIME_BITS'd959819657, `RNS_PRIME_BITS'd852525655},
    '{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd487660555, `RNS_PRIME_BITS'd1061893582, `RNS_PRIME_BITS'd1972644058, `RNS_PRIME_BITS'd812108973, `RNS_PRIME_BITS'd1827722725, `RNS_PRIME_BITS'd285697904, `RNS_PRIME_BITS'd754991627, `RNS_PRIME_BITS'd69473664, `RNS_PRIME_BITS'd1068745859, `RNS_PRIME_BITS'd877540689},
    '{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd1516766091, `RNS_PRIME_BITS'd1468304672, `RNS_PRIME_BITS'd792042504, `RNS_PRIME_BITS'd665252307, `RNS_PRIME_BITS'd1182398267, `RNS_PRIME_BITS'd1478596903, `RNS_PRIME_BITS'd1625334052, `RNS_PRIME_BITS'd1204101513, `RNS_PRIME_BITS'd1517514452, `RNS_PRIME_BITS'd1852392826},
    '{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd235675091, `RNS_PRIME_BITS'd1215871282, `RNS_PRIME_BITS'd1745394775, `RNS_PRIME_BITS'd547832513, `RNS_PRIME_BITS'd832031840, `RNS_PRIME_BITS'd1084796080, `RNS_PRIME_BITS'd1494828160, `RNS_PRIME_BITS'd917052292, `RNS_PRIME_BITS'd1092506897, `RNS_PRIME_BITS'd1715992980},
    '{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd1277622228, `RNS_PRIME_BITS'd687833643, `RNS_PRIME_BITS'd126756375, `RNS_PRIME_BITS'd765208504, `RNS_PRIME_BITS'd1634973533, `RNS_PRIME_BITS'd114865935, `RNS_PRIME_BITS'd491511062, `RNS_PRIME_BITS'd1938597003, `RNS_PRIME_BITS'd715389181, `RNS_PRIME_BITS'd1443341153},
    '{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd1825586477, `RNS_PRIME_BITS'd1396430759, `RNS_PRIME_BITS'd1303407128, `RNS_PRIME_BITS'd1445475149, `RNS_PRIME_BITS'd424619735, `RNS_PRIME_BITS'd41354298, `RNS_PRIME_BITS'd1409837468, `RNS_PRIME_BITS'd278181591, `RNS_PRIME_BITS'd1819301706, `RNS_PRIME_BITS'd1848035921},
    '{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd1904686822, `RNS_PRIME_BITS'd1106318626, `RNS_PRIME_BITS'd644769538, `RNS_PRIME_BITS'd923417179, `RNS_PRIME_BITS'd1061536840, `RNS_PRIME_BITS'd206347908, `RNS_PRIME_BITS'd960907922, `RNS_PRIME_BITS'd2014200918, `RNS_PRIME_BITS'd1799695897, `RNS_PRIME_BITS'd184868460},
    '{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd1660605546, `RNS_PRIME_BITS'd1932790523, `RNS_PRIME_BITS'd107468360, `RNS_PRIME_BITS'd1475935526, `RNS_PRIME_BITS'd2137031813, `RNS_PRIME_BITS'd1842075581, `RNS_PRIME_BITS'd1534159273, `RNS_PRIME_BITS'd1414891420, `RNS_PRIME_BITS'd114674984, `RNS_PRIME_BITS'd422161172},
    '{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd1467716298, `RNS_PRIME_BITS'd1845758024, `RNS_PRIME_BITS'd2027318364, `RNS_PRIME_BITS'd1497830248, `RNS_PRIME_BITS'd1322321168, `RNS_PRIME_BITS'd1937021108, `RNS_PRIME_BITS'd58754948, `RNS_PRIME_BITS'd2075407172, `RNS_PRIME_BITS'd983943721, `RNS_PRIME_BITS'd2147117881},
    '{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd2014655720, `RNS_PRIME_BITS'd1862208197, `RNS_PRIME_BITS'd1311559924, `RNS_PRIME_BITS'd1955877019, `RNS_PRIME_BITS'd2076220394, `RNS_PRIME_BITS'd257564127, `RNS_PRIME_BITS'd565055248, `RNS_PRIME_BITS'd1143569118, `RNS_PRIME_BITS'd791472279, `RNS_PRIME_BITS'd927992919},
    '{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd1680150016, `RNS_PRIME_BITS'd1828982382, `RNS_PRIME_BITS'd250397076, `RNS_PRIME_BITS'd767075907, `RNS_PRIME_BITS'd1216694894, `RNS_PRIME_BITS'd1666228359, `RNS_PRIME_BITS'd1911095743, `RNS_PRIME_BITS'd947926127, `RNS_PRIME_BITS'd69398065, `RNS_PRIME_BITS'd147306452},
    '{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd929720665, `RNS_PRIME_BITS'd1370616561, `RNS_PRIME_BITS'd1312952281, `RNS_PRIME_BITS'd1642055929, `RNS_PRIME_BITS'd1027913888, `RNS_PRIME_BITS'd1836041565, `RNS_PRIME_BITS'd812388307, `RNS_PRIME_BITS'd1235506155, `RNS_PRIME_BITS'd1868402086, `RNS_PRIME_BITS'd197841319},
    '{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd828673995, `RNS_PRIME_BITS'd575270028, `RNS_PRIME_BITS'd620510798, `RNS_PRIME_BITS'd308787199, `RNS_PRIME_BITS'd1057096300, `RNS_PRIME_BITS'd61639648, `RNS_PRIME_BITS'd1980586176, `RNS_PRIME_BITS'd2144543143, `RNS_PRIME_BITS'd1035521899, `RNS_PRIME_BITS'd1481261841},
    '{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd1869944373, `RNS_PRIME_BITS'd1813643879, `RNS_PRIME_BITS'd1870421688, `RNS_PRIME_BITS'd1548197755, `RNS_PRIME_BITS'd1032972630, `RNS_PRIME_BITS'd1961780163, `RNS_PRIME_BITS'd206032257, `RNS_PRIME_BITS'd341345352, `RNS_PRIME_BITS'd1296559053, `RNS_PRIME_BITS'd1100192790},
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1671046886, `RNS_PRIME_BITS'd779176347, `RNS_PRIME_BITS'd395545305, `RNS_PRIME_BITS'd548519104, `RNS_PRIME_BITS'd1521713106, `RNS_PRIME_BITS'd1778166872, `RNS_PRIME_BITS'd1992360836, `RNS_PRIME_BITS'd307943512, `RNS_PRIME_BITS'd1858486778, `RNS_PRIME_BITS'd1217376535},
    '{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd77607433, `RNS_PRIME_BITS'd445781670, `RNS_PRIME_BITS'd362973800, `RNS_PRIME_BITS'd2135267821, `RNS_PRIME_BITS'd762068841, `RNS_PRIME_BITS'd381804377, `RNS_PRIME_BITS'd1356500139, `RNS_PRIME_BITS'd1620634429, `RNS_PRIME_BITS'd846861628, `RNS_PRIME_BITS'd106730909},
    '{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd322709120, `RNS_PRIME_BITS'd834254757, `RNS_PRIME_BITS'd393772305, `RNS_PRIME_BITS'd633431033, `RNS_PRIME_BITS'd1242279121, `RNS_PRIME_BITS'd583416946, `RNS_PRIME_BITS'd609475388, `RNS_PRIME_BITS'd903262245, `RNS_PRIME_BITS'd756641082, `RNS_PRIME_BITS'd236176371},
    '{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd448215137, `RNS_PRIME_BITS'd901976536, `RNS_PRIME_BITS'd445651178, `RNS_PRIME_BITS'd173840560, `RNS_PRIME_BITS'd378485855, `RNS_PRIME_BITS'd1170893215, `RNS_PRIME_BITS'd1404566493, `RNS_PRIME_BITS'd1110642524, `RNS_PRIME_BITS'd366040601, `RNS_PRIME_BITS'd357099177},
    '{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd2067638453, `RNS_PRIME_BITS'd1373132689, `RNS_PRIME_BITS'd773754097, `RNS_PRIME_BITS'd1816808974, `RNS_PRIME_BITS'd717957840, `RNS_PRIME_BITS'd1775229345, `RNS_PRIME_BITS'd333239654, `RNS_PRIME_BITS'd199427305, `RNS_PRIME_BITS'd1605368013, `RNS_PRIME_BITS'd946081369},
    '{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd762782950, `RNS_PRIME_BITS'd1381901223, `RNS_PRIME_BITS'd786873016, `RNS_PRIME_BITS'd451947566, `RNS_PRIME_BITS'd71222797, `RNS_PRIME_BITS'd1750410703, `RNS_PRIME_BITS'd561271880, `RNS_PRIME_BITS'd402400139, `RNS_PRIME_BITS'd822622409, `RNS_PRIME_BITS'd1215563929},
    '{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd1894558169, `RNS_PRIME_BITS'd1252004129, `RNS_PRIME_BITS'd116503006, `RNS_PRIME_BITS'd752064863, `RNS_PRIME_BITS'd218438491, `RNS_PRIME_BITS'd603153407, `RNS_PRIME_BITS'd1408479531, `RNS_PRIME_BITS'd814442837, `RNS_PRIME_BITS'd1190173409, `RNS_PRIME_BITS'd2137012790},
    '{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1366303369, `RNS_PRIME_BITS'd9501924, `RNS_PRIME_BITS'd1040884399, `RNS_PRIME_BITS'd402384571, `RNS_PRIME_BITS'd1181165213, `RNS_PRIME_BITS'd1573770178, `RNS_PRIME_BITS'd1405940624, `RNS_PRIME_BITS'd1024760168, `RNS_PRIME_BITS'd1506088651, `RNS_PRIME_BITS'd1013324149},
    '{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd1144638401, `RNS_PRIME_BITS'd3893692, `RNS_PRIME_BITS'd1435611144, `RNS_PRIME_BITS'd554819808, `RNS_PRIME_BITS'd1532223950, `RNS_PRIME_BITS'd594106318, `RNS_PRIME_BITS'd772678882, `RNS_PRIME_BITS'd305693585, `RNS_PRIME_BITS'd2109818209, `RNS_PRIME_BITS'd980397734},
    '{`RNS_PRIME_BITS'd219, `RNS_PRIME_BITS'd710389119, `RNS_PRIME_BITS'd381253997, `RNS_PRIME_BITS'd930727903, `RNS_PRIME_BITS'd1386770720, `RNS_PRIME_BITS'd891839277, `RNS_PRIME_BITS'd137013315, `RNS_PRIME_BITS'd2077681754, `RNS_PRIME_BITS'd146278937, `RNS_PRIME_BITS'd883007174, `RNS_PRIME_BITS'd152000087},
    '{`RNS_PRIME_BITS'd165, `RNS_PRIME_BITS'd682581400, `RNS_PRIME_BITS'd1455981910, `RNS_PRIME_BITS'd878917060, `RNS_PRIME_BITS'd2041288751, `RNS_PRIME_BITS'd255425535, `RNS_PRIME_BITS'd423747580, `RNS_PRIME_BITS'd1624241031, `RNS_PRIME_BITS'd163998385, `RNS_PRIME_BITS'd1049135090, `RNS_PRIME_BITS'd252484763},
    '{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1397784951, `RNS_PRIME_BITS'd1865708240, `RNS_PRIME_BITS'd2003438866, `RNS_PRIME_BITS'd1733411078, `RNS_PRIME_BITS'd1002091085, `RNS_PRIME_BITS'd1221828305, `RNS_PRIME_BITS'd1999633365, `RNS_PRIME_BITS'd876370933, `RNS_PRIME_BITS'd1885910635, `RNS_PRIME_BITS'd2095966213},
    '{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd1384564752, `RNS_PRIME_BITS'd433472788, `RNS_PRIME_BITS'd665425110, `RNS_PRIME_BITS'd1773817788, `RNS_PRIME_BITS'd213524890, `RNS_PRIME_BITS'd1659723709, `RNS_PRIME_BITS'd1906464361, `RNS_PRIME_BITS'd1552802447, `RNS_PRIME_BITS'd2049845174, `RNS_PRIME_BITS'd1300791096},
    '{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd338600753, `RNS_PRIME_BITS'd1538317438, `RNS_PRIME_BITS'd1105809867, `RNS_PRIME_BITS'd819333801, `RNS_PRIME_BITS'd441715862, `RNS_PRIME_BITS'd1213047921, `RNS_PRIME_BITS'd1804074273, `RNS_PRIME_BITS'd549432341, `RNS_PRIME_BITS'd1371046953, `RNS_PRIME_BITS'd1519781316},
    '{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd2129008001, `RNS_PRIME_BITS'd1965939120, `RNS_PRIME_BITS'd1344460707, `RNS_PRIME_BITS'd1017466165, `RNS_PRIME_BITS'd540703789, `RNS_PRIME_BITS'd615494018, `RNS_PRIME_BITS'd590648200, `RNS_PRIME_BITS'd1184685854, `RNS_PRIME_BITS'd1020954333, `RNS_PRIME_BITS'd544490801},
    '{`RNS_PRIME_BITS'd209, `RNS_PRIME_BITS'd1439719799, `RNS_PRIME_BITS'd557730061, `RNS_PRIME_BITS'd163664946, `RNS_PRIME_BITS'd2060177819, `RNS_PRIME_BITS'd1658964647, `RNS_PRIME_BITS'd102829226, `RNS_PRIME_BITS'd23132681, `RNS_PRIME_BITS'd842827861, `RNS_PRIME_BITS'd67300044, `RNS_PRIME_BITS'd1916779228},
    '{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd216832388, `RNS_PRIME_BITS'd1499638702, `RNS_PRIME_BITS'd215052704, `RNS_PRIME_BITS'd889904893, `RNS_PRIME_BITS'd992089543, `RNS_PRIME_BITS'd1968596455, `RNS_PRIME_BITS'd1877331516, `RNS_PRIME_BITS'd1711973714, `RNS_PRIME_BITS'd1056600617, `RNS_PRIME_BITS'd1040737733},
    '{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd1064824235, `RNS_PRIME_BITS'd987830523, `RNS_PRIME_BITS'd827448682, `RNS_PRIME_BITS'd1881048101, `RNS_PRIME_BITS'd77131150, `RNS_PRIME_BITS'd1431760059, `RNS_PRIME_BITS'd671022630, `RNS_PRIME_BITS'd1632059779, `RNS_PRIME_BITS'd147984288, `RNS_PRIME_BITS'd444699212},
    '{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd446909929, `RNS_PRIME_BITS'd1145656905, `RNS_PRIME_BITS'd87751062, `RNS_PRIME_BITS'd651823414, `RNS_PRIME_BITS'd2111085037, `RNS_PRIME_BITS'd1283873057, `RNS_PRIME_BITS'd435908200, `RNS_PRIME_BITS'd989349162, `RNS_PRIME_BITS'd1066794502, `RNS_PRIME_BITS'd751065570},
    '{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd2035000636, `RNS_PRIME_BITS'd1299571809, `RNS_PRIME_BITS'd397159397, `RNS_PRIME_BITS'd1149497610, `RNS_PRIME_BITS'd285868357, `RNS_PRIME_BITS'd860170220, `RNS_PRIME_BITS'd957433122, `RNS_PRIME_BITS'd1648166161, `RNS_PRIME_BITS'd1850235833, `RNS_PRIME_BITS'd1790613488},
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1013199338, `RNS_PRIME_BITS'd1968587998, `RNS_PRIME_BITS'd1289695665, `RNS_PRIME_BITS'd296590121, `RNS_PRIME_BITS'd280092226, `RNS_PRIME_BITS'd2063421943, `RNS_PRIME_BITS'd901372286, `RNS_PRIME_BITS'd737217449, `RNS_PRIME_BITS'd1532531378, `RNS_PRIME_BITS'd1550494478},
    '{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd299380480, `RNS_PRIME_BITS'd255743251, `RNS_PRIME_BITS'd1788013446, `RNS_PRIME_BITS'd2049595553, `RNS_PRIME_BITS'd253819890, `RNS_PRIME_BITS'd162154740, `RNS_PRIME_BITS'd928213509, `RNS_PRIME_BITS'd718679450, `RNS_PRIME_BITS'd671227245, `RNS_PRIME_BITS'd572242555},
    '{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd667783287, `RNS_PRIME_BITS'd794056254, `RNS_PRIME_BITS'd39422024, `RNS_PRIME_BITS'd170203145, `RNS_PRIME_BITS'd972447735, `RNS_PRIME_BITS'd1332479475, `RNS_PRIME_BITS'd714672611, `RNS_PRIME_BITS'd2109603880, `RNS_PRIME_BITS'd571950693, `RNS_PRIME_BITS'd762736245},
    '{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd1115696555, `RNS_PRIME_BITS'd1538380880, `RNS_PRIME_BITS'd1548856345, `RNS_PRIME_BITS'd1472321400, `RNS_PRIME_BITS'd1043517755, `RNS_PRIME_BITS'd922417491, `RNS_PRIME_BITS'd2049492523, `RNS_PRIME_BITS'd212262096, `RNS_PRIME_BITS'd619627638, `RNS_PRIME_BITS'd1503925676},
    '{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd1777896165, `RNS_PRIME_BITS'd1394135005, `RNS_PRIME_BITS'd1526298610, `RNS_PRIME_BITS'd1881386209, `RNS_PRIME_BITS'd996757604, `RNS_PRIME_BITS'd1031386265, `RNS_PRIME_BITS'd1905368146, `RNS_PRIME_BITS'd130410828, `RNS_PRIME_BITS'd717318262, `RNS_PRIME_BITS'd1885797622},
    '{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd1489514692, `RNS_PRIME_BITS'd399680613, `RNS_PRIME_BITS'd1884286346, `RNS_PRIME_BITS'd79271719, `RNS_PRIME_BITS'd1697376542, `RNS_PRIME_BITS'd973747397, `RNS_PRIME_BITS'd540796709, `RNS_PRIME_BITS'd2020879262, `RNS_PRIME_BITS'd1194089328, `RNS_PRIME_BITS'd673980632},
    '{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd961661966, `RNS_PRIME_BITS'd1775541313, `RNS_PRIME_BITS'd243665668, `RNS_PRIME_BITS'd845308960, `RNS_PRIME_BITS'd1018410470, `RNS_PRIME_BITS'd1792340588, `RNS_PRIME_BITS'd2076560098, `RNS_PRIME_BITS'd894044508, `RNS_PRIME_BITS'd740049617, `RNS_PRIME_BITS'd442752118},
    '{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd490495528, `RNS_PRIME_BITS'd218892080, `RNS_PRIME_BITS'd258539907, `RNS_PRIME_BITS'd1967225852, `RNS_PRIME_BITS'd657983768, `RNS_PRIME_BITS'd948953814, `RNS_PRIME_BITS'd636783003, `RNS_PRIME_BITS'd729293999, `RNS_PRIME_BITS'd814288155, `RNS_PRIME_BITS'd93362422},
    '{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd1412279211, `RNS_PRIME_BITS'd40804773, `RNS_PRIME_BITS'd405570514, `RNS_PRIME_BITS'd1438162702, `RNS_PRIME_BITS'd1946144078, `RNS_PRIME_BITS'd330336588, `RNS_PRIME_BITS'd1397243825, `RNS_PRIME_BITS'd1449491717, `RNS_PRIME_BITS'd1477538017, `RNS_PRIME_BITS'd1177794342},
    '{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd1110789405, `RNS_PRIME_BITS'd626528868, `RNS_PRIME_BITS'd881138703, `RNS_PRIME_BITS'd1933195299, `RNS_PRIME_BITS'd1114586919, `RNS_PRIME_BITS'd821409919, `RNS_PRIME_BITS'd130646675, `RNS_PRIME_BITS'd1873235257, `RNS_PRIME_BITS'd1690386107, `RNS_PRIME_BITS'd721418499},
    '{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd1484266757, `RNS_PRIME_BITS'd1300731878, `RNS_PRIME_BITS'd1409114395, `RNS_PRIME_BITS'd1846628098, `RNS_PRIME_BITS'd980139663, `RNS_PRIME_BITS'd703773412, `RNS_PRIME_BITS'd1197908194, `RNS_PRIME_BITS'd626823517, `RNS_PRIME_BITS'd1621578307, `RNS_PRIME_BITS'd635217709},
    '{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd734332099, `RNS_PRIME_BITS'd498345152, `RNS_PRIME_BITS'd692737758, `RNS_PRIME_BITS'd1662562743, `RNS_PRIME_BITS'd1541319866, `RNS_PRIME_BITS'd1270899383, `RNS_PRIME_BITS'd1458093008, `RNS_PRIME_BITS'd760536533, `RNS_PRIME_BITS'd1507237810, `RNS_PRIME_BITS'd1939598861},
    '{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd2089344066, `RNS_PRIME_BITS'd544473085, `RNS_PRIME_BITS'd1714517841, `RNS_PRIME_BITS'd1913047875, `RNS_PRIME_BITS'd625018383, `RNS_PRIME_BITS'd1267544990, `RNS_PRIME_BITS'd638371721, `RNS_PRIME_BITS'd1705055400, `RNS_PRIME_BITS'd1433120257, `RNS_PRIME_BITS'd525740258},
    '{`RNS_PRIME_BITS'd10, `RNS_PRIME_BITS'd414159494, `RNS_PRIME_BITS'd163452829, `RNS_PRIME_BITS'd2111205207, `RNS_PRIME_BITS'd1605954173, `RNS_PRIME_BITS'd976805569, `RNS_PRIME_BITS'd2088726651, `RNS_PRIME_BITS'd935565441, `RNS_PRIME_BITS'd80201478, `RNS_PRIME_BITS'd397089621, `RNS_PRIME_BITS'd783202583},
    '{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd1147595380, `RNS_PRIME_BITS'd1641914833, `RNS_PRIME_BITS'd1574531044, `RNS_PRIME_BITS'd21766817, `RNS_PRIME_BITS'd1653584508, `RNS_PRIME_BITS'd1868863705, `RNS_PRIME_BITS'd1930662801, `RNS_PRIME_BITS'd782387793, `RNS_PRIME_BITS'd370535898, `RNS_PRIME_BITS'd1969474147},
    '{`RNS_PRIME_BITS'd110, `RNS_PRIME_BITS'd338759259, `RNS_PRIME_BITS'd132866527, `RNS_PRIME_BITS'd462337302, `RNS_PRIME_BITS'd1810257211, `RNS_PRIME_BITS'd271485432, `RNS_PRIME_BITS'd2092074032, `RNS_PRIME_BITS'd1225657871, `RNS_PRIME_BITS'd1816845920, `RNS_PRIME_BITS'd241185360, `RNS_PRIME_BITS'd845414760},
    '{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd1747421548, `RNS_PRIME_BITS'd4671678, `RNS_PRIME_BITS'd1007692149, `RNS_PRIME_BITS'd1622924542, `RNS_PRIME_BITS'd1657536354, `RNS_PRIME_BITS'd1511478571, `RNS_PRIME_BITS'd731731277, `RNS_PRIME_BITS'd767316846, `RNS_PRIME_BITS'd1078196739, `RNS_PRIME_BITS'd1471576852},
    '{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd1786397361, `RNS_PRIME_BITS'd1613071122, `RNS_PRIME_BITS'd2113126473, `RNS_PRIME_BITS'd1684716348, `RNS_PRIME_BITS'd144713126, `RNS_PRIME_BITS'd1880867112, `RNS_PRIME_BITS'd538142292, `RNS_PRIME_BITS'd1997060930, `RNS_PRIME_BITS'd1552885288, `RNS_PRIME_BITS'd1889412258}
};


const rns_residue_t B1__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd1112177129, `RNS_PRIME_BITS'd533724018, `RNS_PRIME_BITS'd177369642, `RNS_PRIME_BITS'd1679005539, `RNS_PRIME_BITS'd53351151, `RNS_PRIME_BITS'd2070494231, `RNS_PRIME_BITS'd1541419757, `RNS_PRIME_BITS'd1696370584, `RNS_PRIME_BITS'd347098394, `RNS_PRIME_BITS'd437246425},
    '{`RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd1073643522, `RNS_PRIME_BITS'd1839593151, `RNS_PRIME_BITS'd1737833868, `RNS_PRIME_BITS'd475564002, `RNS_PRIME_BITS'd1170319951, `RNS_PRIME_BITS'd1652591676, `RNS_PRIME_BITS'd1893033483, `RNS_PRIME_BITS'd1289139607, `RNS_PRIME_BITS'd1822810014, `RNS_PRIME_BITS'd901509048},
    '{`RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd1573781464, `RNS_PRIME_BITS'd993476670, `RNS_PRIME_BITS'd1507418709, `RNS_PRIME_BITS'd874189346, `RNS_PRIME_BITS'd692173684, `RNS_PRIME_BITS'd1932035896, `RNS_PRIME_BITS'd102459851, `RNS_PRIME_BITS'd954571406, `RNS_PRIME_BITS'd326083751, `RNS_PRIME_BITS'd1858900646},
    '{`RNS_PRIME_BITS'd40, `RNS_PRIME_BITS'd642013974, `RNS_PRIME_BITS'd330177291, `RNS_PRIME_BITS'd1879332416, `RNS_PRIME_BITS'd427739881, `RNS_PRIME_BITS'd26936754, `RNS_PRIME_BITS'd532533065, `RNS_PRIME_BITS'd238101500, `RNS_PRIME_BITS'd353341552, `RNS_PRIME_BITS'd1979250593, `RNS_PRIME_BITS'd1650878797},
    '{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd1535568653, `RNS_PRIME_BITS'd1348127996, `RNS_PRIME_BITS'd1184988661, `RNS_PRIME_BITS'd775725997, `RNS_PRIME_BITS'd1284421049, `RNS_PRIME_BITS'd1875436923, `RNS_PRIME_BITS'd555592030, `RNS_PRIME_BITS'd1809645726, `RNS_PRIME_BITS'd421487265, `RNS_PRIME_BITS'd1836811101},
    '{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd1805432572, `RNS_PRIME_BITS'd1479444956, `RNS_PRIME_BITS'd244255772, `RNS_PRIME_BITS'd1224792621, `RNS_PRIME_BITS'd319799473, `RNS_PRIME_BITS'd347843552, `RNS_PRIME_BITS'd36778632, `RNS_PRIME_BITS'd675486343, `RNS_PRIME_BITS'd2009285989, `RNS_PRIME_BITS'd294120590},
    '{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1986164302, `RNS_PRIME_BITS'd1598529123, `RNS_PRIME_BITS'd1436650056, `RNS_PRIME_BITS'd1643346754, `RNS_PRIME_BITS'd272751409, `RNS_PRIME_BITS'd2007774725, `RNS_PRIME_BITS'd709297183, `RNS_PRIME_BITS'd75598114, `RNS_PRIME_BITS'd559874540, `RNS_PRIME_BITS'd2069463412},
    '{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd1573748397, `RNS_PRIME_BITS'd454327866, `RNS_PRIME_BITS'd1498198573, `RNS_PRIME_BITS'd2111692288, `RNS_PRIME_BITS'd49349786, `RNS_PRIME_BITS'd1863696370, `RNS_PRIME_BITS'd1862307613, `RNS_PRIME_BITS'd695707078, `RNS_PRIME_BITS'd1806252202, `RNS_PRIME_BITS'd285885355},
    '{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd793712967, `RNS_PRIME_BITS'd1379276324, `RNS_PRIME_BITS'd940594249, `RNS_PRIME_BITS'd251432030, `RNS_PRIME_BITS'd1054277902, `RNS_PRIME_BITS'd1259679508, `RNS_PRIME_BITS'd1875681121, `RNS_PRIME_BITS'd94997646, `RNS_PRIME_BITS'd1179282861, `RNS_PRIME_BITS'd1651078169},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1175247393, `RNS_PRIME_BITS'd1859984809, `RNS_PRIME_BITS'd1570158002, `RNS_PRIME_BITS'd686201950, `RNS_PRIME_BITS'd1310180575, `RNS_PRIME_BITS'd224171677, `RNS_PRIME_BITS'd358778910, `RNS_PRIME_BITS'd1044836134, `RNS_PRIME_BITS'd1536609293, `RNS_PRIME_BITS'd996445963},
    '{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd1209786132, `RNS_PRIME_BITS'd120134476, `RNS_PRIME_BITS'd542613024, `RNS_PRIME_BITS'd1303774552, `RNS_PRIME_BITS'd1945101819, `RNS_PRIME_BITS'd1838674286, `RNS_PRIME_BITS'd2099921013, `RNS_PRIME_BITS'd1995139140, `RNS_PRIME_BITS'd216989534, `RNS_PRIME_BITS'd1052103703},
    '{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd323465263, `RNS_PRIME_BITS'd1919920336, `RNS_PRIME_BITS'd2120776927, `RNS_PRIME_BITS'd1636300436, `RNS_PRIME_BITS'd1539610205, `RNS_PRIME_BITS'd155259357, `RNS_PRIME_BITS'd1954766997, `RNS_PRIME_BITS'd585577790, `RNS_PRIME_BITS'd1447080486, `RNS_PRIME_BITS'd623930340},
    '{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd1317357696, `RNS_PRIME_BITS'd563472138, `RNS_PRIME_BITS'd1848835296, `RNS_PRIME_BITS'd1030568412, `RNS_PRIME_BITS'd473560242, `RNS_PRIME_BITS'd303622602, `RNS_PRIME_BITS'd258042911, `RNS_PRIME_BITS'd1350930064, `RNS_PRIME_BITS'd1206935249, `RNS_PRIME_BITS'd2026007438},
    '{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd273472676, `RNS_PRIME_BITS'd1009731306, `RNS_PRIME_BITS'd1449642614, `RNS_PRIME_BITS'd552032419, `RNS_PRIME_BITS'd1095771470, `RNS_PRIME_BITS'd1077074841, `RNS_PRIME_BITS'd2009540477, `RNS_PRIME_BITS'd1904124804, `RNS_PRIME_BITS'd1728187142, `RNS_PRIME_BITS'd39381268},
    '{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd114973466, `RNS_PRIME_BITS'd1032654110, `RNS_PRIME_BITS'd424623646, `RNS_PRIME_BITS'd622386704, `RNS_PRIME_BITS'd958463837, `RNS_PRIME_BITS'd2083997396, `RNS_PRIME_BITS'd463044865, `RNS_PRIME_BITS'd1928399822, `RNS_PRIME_BITS'd1147380492, `RNS_PRIME_BITS'd1306913883},
    '{`RNS_PRIME_BITS'd127, `RNS_PRIME_BITS'd205335062, `RNS_PRIME_BITS'd1886108378, `RNS_PRIME_BITS'd417507716, `RNS_PRIME_BITS'd1311297208, `RNS_PRIME_BITS'd1761787573, `RNS_PRIME_BITS'd733919294, `RNS_PRIME_BITS'd379871042, `RNS_PRIME_BITS'd1672289110, `RNS_PRIME_BITS'd2033261300, `RNS_PRIME_BITS'd470497662},
    '{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd929474099, `RNS_PRIME_BITS'd931895367, `RNS_PRIME_BITS'd1135264550, `RNS_PRIME_BITS'd904652825, `RNS_PRIME_BITS'd26041371, `RNS_PRIME_BITS'd1282426128, `RNS_PRIME_BITS'd325859244, `RNS_PRIME_BITS'd285135055, `RNS_PRIME_BITS'd1076641534, `RNS_PRIME_BITS'd781758218},
    '{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd2087640943, `RNS_PRIME_BITS'd111135999, `RNS_PRIME_BITS'd603708949, `RNS_PRIME_BITS'd1834610488, `RNS_PRIME_BITS'd1555370594, `RNS_PRIME_BITS'd2081115710, `RNS_PRIME_BITS'd1997540534, `RNS_PRIME_BITS'd1116957688, `RNS_PRIME_BITS'd41882368, `RNS_PRIME_BITS'd829777403},
    '{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd1137914064, `RNS_PRIME_BITS'd1836344921, `RNS_PRIME_BITS'd520131278, `RNS_PRIME_BITS'd38364964, `RNS_PRIME_BITS'd1536109204, `RNS_PRIME_BITS'd1684360183, `RNS_PRIME_BITS'd905999784, `RNS_PRIME_BITS'd713215541, `RNS_PRIME_BITS'd474109682, `RNS_PRIME_BITS'd37534420},
    '{`RNS_PRIME_BITS'd254, `RNS_PRIME_BITS'd50724854, `RNS_PRIME_BITS'd441216682, `RNS_PRIME_BITS'd1558450071, `RNS_PRIME_BITS'd175251213, `RNS_PRIME_BITS'd1427316831, `RNS_PRIME_BITS'd1325475735, `RNS_PRIME_BITS'd1883296115, `RNS_PRIME_BITS'd972722944, `RNS_PRIME_BITS'd591159602, `RNS_PRIME_BITS'd1257059938},
    '{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd1790526299, `RNS_PRIME_BITS'd1142469266, `RNS_PRIME_BITS'd846814023, `RNS_PRIME_BITS'd1632341828, `RNS_PRIME_BITS'd686687228, `RNS_PRIME_BITS'd1030300001, `RNS_PRIME_BITS'd885556596, `RNS_PRIME_BITS'd300196478, `RNS_PRIME_BITS'd2118400297, `RNS_PRIME_BITS'd2120870941},
    '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd274699930, `RNS_PRIME_BITS'd251379313, `RNS_PRIME_BITS'd1526905374, `RNS_PRIME_BITS'd122336816, `RNS_PRIME_BITS'd341917250, `RNS_PRIME_BITS'd1485190407, `RNS_PRIME_BITS'd1444780686, `RNS_PRIME_BITS'd1826772569, `RNS_PRIME_BITS'd280136862, `RNS_PRIME_BITS'd99978015},
    '{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd856480772, `RNS_PRIME_BITS'd1599804981, `RNS_PRIME_BITS'd2118686352, `RNS_PRIME_BITS'd2092037920, `RNS_PRIME_BITS'd747563730, `RNS_PRIME_BITS'd2060261769, `RNS_PRIME_BITS'd1561048655, `RNS_PRIME_BITS'd1061630524, `RNS_PRIME_BITS'd1455980167, `RNS_PRIME_BITS'd242505757},
    '{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd1974415341, `RNS_PRIME_BITS'd119315056, `RNS_PRIME_BITS'd1564842323, `RNS_PRIME_BITS'd1660438749, `RNS_PRIME_BITS'd1550063706, `RNS_PRIME_BITS'd717930396, `RNS_PRIME_BITS'd1211259340, `RNS_PRIME_BITS'd1241714252, `RNS_PRIME_BITS'd793254048, `RNS_PRIME_BITS'd846536775},
    '{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd143359173, `RNS_PRIME_BITS'd172540774, `RNS_PRIME_BITS'd932916068, `RNS_PRIME_BITS'd1922634531, `RNS_PRIME_BITS'd1868506357, `RNS_PRIME_BITS'd714680179, `RNS_PRIME_BITS'd1074790157, `RNS_PRIME_BITS'd1345953698, `RNS_PRIME_BITS'd2128692625, `RNS_PRIME_BITS'd202642545},
    '{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd1117142210, `RNS_PRIME_BITS'd1679150616, `RNS_PRIME_BITS'd528529137, `RNS_PRIME_BITS'd1873055888, `RNS_PRIME_BITS'd2015238493, `RNS_PRIME_BITS'd718828362, `RNS_PRIME_BITS'd2144090113, `RNS_PRIME_BITS'd676470118, `RNS_PRIME_BITS'd96294373, `RNS_PRIME_BITS'd1772680642},
    '{`RNS_PRIME_BITS'd127, `RNS_PRIME_BITS'd996309165, `RNS_PRIME_BITS'd1207918232, `RNS_PRIME_BITS'd807082959, `RNS_PRIME_BITS'd1936000263, `RNS_PRIME_BITS'd751961263, `RNS_PRIME_BITS'd1436729800, `RNS_PRIME_BITS'd1193790209, `RNS_PRIME_BITS'd2037821185, `RNS_PRIME_BITS'd1037098591, `RNS_PRIME_BITS'd1288545473},
    '{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd833129398, `RNS_PRIME_BITS'd1902828236, `RNS_PRIME_BITS'd930672877, `RNS_PRIME_BITS'd228521520, `RNS_PRIME_BITS'd922443347, `RNS_PRIME_BITS'd1348733276, `RNS_PRIME_BITS'd2075809, `RNS_PRIME_BITS'd1161009867, `RNS_PRIME_BITS'd1292162686, `RNS_PRIME_BITS'd12766120},
    '{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd790372, `RNS_PRIME_BITS'd81104610, `RNS_PRIME_BITS'd1539322725, `RNS_PRIME_BITS'd707502649, `RNS_PRIME_BITS'd575965510, `RNS_PRIME_BITS'd283699902, `RNS_PRIME_BITS'd347711999, `RNS_PRIME_BITS'd1982566773, `RNS_PRIME_BITS'd968607687, `RNS_PRIME_BITS'd205361198},
    '{`RNS_PRIME_BITS'd227, `RNS_PRIME_BITS'd1697214269, `RNS_PRIME_BITS'd2070533898, `RNS_PRIME_BITS'd1249720436, `RNS_PRIME_BITS'd1338706744, `RNS_PRIME_BITS'd1732282581, `RNS_PRIME_BITS'd250645440, `RNS_PRIME_BITS'd2059198497, `RNS_PRIME_BITS'd566771231, `RNS_PRIME_BITS'd1647576202, `RNS_PRIME_BITS'd1653833293},
    '{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd629085881, `RNS_PRIME_BITS'd617284009, `RNS_PRIME_BITS'd1259963447, `RNS_PRIME_BITS'd479018809, `RNS_PRIME_BITS'd57176881, `RNS_PRIME_BITS'd406981233, `RNS_PRIME_BITS'd299561556, `RNS_PRIME_BITS'd1919910668, `RNS_PRIME_BITS'd837949126, `RNS_PRIME_BITS'd392964044},
    '{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd1155221625, `RNS_PRIME_BITS'd1115962718, `RNS_PRIME_BITS'd1107701069, `RNS_PRIME_BITS'd1884712943, `RNS_PRIME_BITS'd1906075553, `RNS_PRIME_BITS'd1485486612, `RNS_PRIME_BITS'd11167576, `RNS_PRIME_BITS'd1120042161, `RNS_PRIME_BITS'd567908485, `RNS_PRIME_BITS'd224547886},
    '{`RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd1965386384, `RNS_PRIME_BITS'd269005161, `RNS_PRIME_BITS'd242053564, `RNS_PRIME_BITS'd610786302, `RNS_PRIME_BITS'd1838563798, `RNS_PRIME_BITS'd1476567249, `RNS_PRIME_BITS'd2059693533, `RNS_PRIME_BITS'd1777827796, `RNS_PRIME_BITS'd670852388, `RNS_PRIME_BITS'd844248888},
    '{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd1134339826, `RNS_PRIME_BITS'd374409069, `RNS_PRIME_BITS'd1712228255, `RNS_PRIME_BITS'd1494014664, `RNS_PRIME_BITS'd1111161830, `RNS_PRIME_BITS'd111038966, `RNS_PRIME_BITS'd2002186540, `RNS_PRIME_BITS'd1207964588, `RNS_PRIME_BITS'd1283198888, `RNS_PRIME_BITS'd307022269},
    '{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd951055158, `RNS_PRIME_BITS'd1324536093, `RNS_PRIME_BITS'd627027284, `RNS_PRIME_BITS'd1306671701, `RNS_PRIME_BITS'd464939954, `RNS_PRIME_BITS'd295729342, `RNS_PRIME_BITS'd828055864, `RNS_PRIME_BITS'd1213152909, `RNS_PRIME_BITS'd1335574470, `RNS_PRIME_BITS'd1376581910},
    '{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd1540780196, `RNS_PRIME_BITS'd587249532, `RNS_PRIME_BITS'd685733135, `RNS_PRIME_BITS'd1621209726, `RNS_PRIME_BITS'd48171582, `RNS_PRIME_BITS'd141561841, `RNS_PRIME_BITS'd1252461035, `RNS_PRIME_BITS'd1787854826, `RNS_PRIME_BITS'd960780260, `RNS_PRIME_BITS'd1444163481},
    '{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1772712583, `RNS_PRIME_BITS'd82039703, `RNS_PRIME_BITS'd348823278, `RNS_PRIME_BITS'd1409838555, `RNS_PRIME_BITS'd1534338606, `RNS_PRIME_BITS'd1532893202, `RNS_PRIME_BITS'd536058282, `RNS_PRIME_BITS'd1312782605, `RNS_PRIME_BITS'd1973604921, `RNS_PRIME_BITS'd702817201},
    '{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd684799169, `RNS_PRIME_BITS'd810617567, `RNS_PRIME_BITS'd1563868315, `RNS_PRIME_BITS'd2132277026, `RNS_PRIME_BITS'd1176205619, `RNS_PRIME_BITS'd1291617213, `RNS_PRIME_BITS'd1838737580, `RNS_PRIME_BITS'd1344807810, `RNS_PRIME_BITS'd205029333, `RNS_PRIME_BITS'd1054039332},
    '{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1957191822, `RNS_PRIME_BITS'd713610746, `RNS_PRIME_BITS'd1022258106, `RNS_PRIME_BITS'd137282309, `RNS_PRIME_BITS'd1747397999, `RNS_PRIME_BITS'd1678452135, `RNS_PRIME_BITS'd1374050501, `RNS_PRIME_BITS'd58494818, `RNS_PRIME_BITS'd1920146035, `RNS_PRIME_BITS'd1030312990},
    '{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd1516519767, `RNS_PRIME_BITS'd153726826, `RNS_PRIME_BITS'd481122877, `RNS_PRIME_BITS'd1653785398, `RNS_PRIME_BITS'd1746494811, `RNS_PRIME_BITS'd1421695236, `RNS_PRIME_BITS'd1121160833, `RNS_PRIME_BITS'd1275308650, `RNS_PRIME_BITS'd1539636806, `RNS_PRIME_BITS'd333468000},
    '{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd10127593, `RNS_PRIME_BITS'd1000689173, `RNS_PRIME_BITS'd313552563, `RNS_PRIME_BITS'd676065904, `RNS_PRIME_BITS'd622357238, `RNS_PRIME_BITS'd949605323, `RNS_PRIME_BITS'd384385278, `RNS_PRIME_BITS'd39249878, `RNS_PRIME_BITS'd1197981333, `RNS_PRIME_BITS'd949137539},
    '{`RNS_PRIME_BITS'd200, `RNS_PRIME_BITS'd337931371, `RNS_PRIME_BITS'd1883587920, `RNS_PRIME_BITS'd2144223167, `RNS_PRIME_BITS'd855614653, `RNS_PRIME_BITS'd1520467348, `RNS_PRIME_BITS'd94829644, `RNS_PRIME_BITS'd1404149427, `RNS_PRIME_BITS'd1447443135, `RNS_PRIME_BITS'd1153651156, `RNS_PRIME_BITS'd1330699208},
    '{`RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd2059688595, `RNS_PRIME_BITS'd1667457803, `RNS_PRIME_BITS'd1704998218, `RNS_PRIME_BITS'd212898690, `RNS_PRIME_BITS'd1283772962, `RNS_PRIME_BITS'd1816058201, `RNS_PRIME_BITS'd1838322638, `RNS_PRIME_BITS'd1715861536, `RNS_PRIME_BITS'd1275659246, `RNS_PRIME_BITS'd420883519},
    '{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd100752789, `RNS_PRIME_BITS'd1003691477, `RNS_PRIME_BITS'd1891578876, `RNS_PRIME_BITS'd17834092, `RNS_PRIME_BITS'd760348902, `RNS_PRIME_BITS'd1518570042, `RNS_PRIME_BITS'd803557866, `RNS_PRIME_BITS'd289166600, `RNS_PRIME_BITS'd1465043887, `RNS_PRIME_BITS'd803412716},
    '{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd1717345786, `RNS_PRIME_BITS'd1366360350, `RNS_PRIME_BITS'd23323037, `RNS_PRIME_BITS'd1158294021, `RNS_PRIME_BITS'd1463842813, `RNS_PRIME_BITS'd618382166, `RNS_PRIME_BITS'd2089062549, `RNS_PRIME_BITS'd323297973, `RNS_PRIME_BITS'd1548543636, `RNS_PRIME_BITS'd984931703},
    '{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd937164560, `RNS_PRIME_BITS'd2051324300, `RNS_PRIME_BITS'd1359881549, `RNS_PRIME_BITS'd1048106073, `RNS_PRIME_BITS'd197283874, `RNS_PRIME_BITS'd1088081971, `RNS_PRIME_BITS'd600312126, `RNS_PRIME_BITS'd860429776, `RNS_PRIME_BITS'd1631863014, `RNS_PRIME_BITS'd873653664},
    '{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd199733383, `RNS_PRIME_BITS'd1229117, `RNS_PRIME_BITS'd581351259, `RNS_PRIME_BITS'd400306786, `RNS_PRIME_BITS'd1275471541, `RNS_PRIME_BITS'd1314617843, `RNS_PRIME_BITS'd871309138, `RNS_PRIME_BITS'd507070489, `RNS_PRIME_BITS'd72930674, `RNS_PRIME_BITS'd264662273},
    '{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd1535323094, `RNS_PRIME_BITS'd2110171527, `RNS_PRIME_BITS'd181617893, `RNS_PRIME_BITS'd1240107990, `RNS_PRIME_BITS'd1760785827, `RNS_PRIME_BITS'd625690953, `RNS_PRIME_BITS'd918847505, `RNS_PRIME_BITS'd1121377264, `RNS_PRIME_BITS'd913794679, `RNS_PRIME_BITS'd176667167},
    '{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd1524898395, `RNS_PRIME_BITS'd328776345, `RNS_PRIME_BITS'd1478926208, `RNS_PRIME_BITS'd638627156, `RNS_PRIME_BITS'd1525155909, `RNS_PRIME_BITS'd190214828, `RNS_PRIME_BITS'd939014540, `RNS_PRIME_BITS'd1370006502, `RNS_PRIME_BITS'd1472770741, `RNS_PRIME_BITS'd1901673831},
    '{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd1977356418, `RNS_PRIME_BITS'd1416042109, `RNS_PRIME_BITS'd1268940097, `RNS_PRIME_BITS'd1599005507, `RNS_PRIME_BITS'd1360518250, `RNS_PRIME_BITS'd1852933214, `RNS_PRIME_BITS'd1845618623, `RNS_PRIME_BITS'd1221987483, `RNS_PRIME_BITS'd1025654897, `RNS_PRIME_BITS'd2022986731},
    '{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd1924168720, `RNS_PRIME_BITS'd1117521150, `RNS_PRIME_BITS'd1349322215, `RNS_PRIME_BITS'd1825385250, `RNS_PRIME_BITS'd722760804, `RNS_PRIME_BITS'd1514640852, `RNS_PRIME_BITS'd713033628, `RNS_PRIME_BITS'd1186258765, `RNS_PRIME_BITS'd2082051840, `RNS_PRIME_BITS'd665342043},
    '{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd1624957880, `RNS_PRIME_BITS'd1323885443, `RNS_PRIME_BITS'd105666160, `RNS_PRIME_BITS'd1300983831, `RNS_PRIME_BITS'd1840544031, `RNS_PRIME_BITS'd1383379924, `RNS_PRIME_BITS'd922984323, `RNS_PRIME_BITS'd19271485, `RNS_PRIME_BITS'd270741063, `RNS_PRIME_BITS'd432310070},
    '{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd1783258658, `RNS_PRIME_BITS'd1233720020, `RNS_PRIME_BITS'd2057058459, `RNS_PRIME_BITS'd932263644, `RNS_PRIME_BITS'd1711607142, `RNS_PRIME_BITS'd922882244, `RNS_PRIME_BITS'd2003002428, `RNS_PRIME_BITS'd1659266436, `RNS_PRIME_BITS'd1540243117, `RNS_PRIME_BITS'd1212675656},
    '{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd767797461, `RNS_PRIME_BITS'd449130899, `RNS_PRIME_BITS'd487780480, `RNS_PRIME_BITS'd912922912, `RNS_PRIME_BITS'd805659669, `RNS_PRIME_BITS'd1076739182, `RNS_PRIME_BITS'd1976663148, `RNS_PRIME_BITS'd102864023, `RNS_PRIME_BITS'd1144022462, `RNS_PRIME_BITS'd570311396},
    '{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd1787518897, `RNS_PRIME_BITS'd2129617489, `RNS_PRIME_BITS'd1795316463, `RNS_PRIME_BITS'd1508132779, `RNS_PRIME_BITS'd910772726, `RNS_PRIME_BITS'd823915451, `RNS_PRIME_BITS'd1567449857, `RNS_PRIME_BITS'd1749834906, `RNS_PRIME_BITS'd1936884195, `RNS_PRIME_BITS'd416712942},
    '{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1880538070, `RNS_PRIME_BITS'd1797055427, `RNS_PRIME_BITS'd1032899401, `RNS_PRIME_BITS'd28386578, `RNS_PRIME_BITS'd933519243, `RNS_PRIME_BITS'd2015643943, `RNS_PRIME_BITS'd587367817, `RNS_PRIME_BITS'd575599096, `RNS_PRIME_BITS'd963794549, `RNS_PRIME_BITS'd322785847},
    '{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1767143483, `RNS_PRIME_BITS'd1171034280, `RNS_PRIME_BITS'd801826114, `RNS_PRIME_BITS'd129903153, `RNS_PRIME_BITS'd1285551012, `RNS_PRIME_BITS'd98640461, `RNS_PRIME_BITS'd1499448649, `RNS_PRIME_BITS'd213863183, `RNS_PRIME_BITS'd990285518, `RNS_PRIME_BITS'd564816725},
    '{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd349263378, `RNS_PRIME_BITS'd1725167867, `RNS_PRIME_BITS'd294977853, `RNS_PRIME_BITS'd1364875384, `RNS_PRIME_BITS'd1630016139, `RNS_PRIME_BITS'd20313273, `RNS_PRIME_BITS'd959416456, `RNS_PRIME_BITS'd1023240651, `RNS_PRIME_BITS'd844469708, `RNS_PRIME_BITS'd756943719},
    '{`RNS_PRIME_BITS'd233, `RNS_PRIME_BITS'd287220864, `RNS_PRIME_BITS'd1433201783, `RNS_PRIME_BITS'd1598528648, `RNS_PRIME_BITS'd1239915840, `RNS_PRIME_BITS'd940797769, `RNS_PRIME_BITS'd922005843, `RNS_PRIME_BITS'd552867908, `RNS_PRIME_BITS'd180967113, `RNS_PRIME_BITS'd1437316834, `RNS_PRIME_BITS'd452718313},
    '{`RNS_PRIME_BITS'd210, `RNS_PRIME_BITS'd1580529677, `RNS_PRIME_BITS'd230279241, `RNS_PRIME_BITS'd743086193, `RNS_PRIME_BITS'd532454818, `RNS_PRIME_BITS'd1607468250, `RNS_PRIME_BITS'd966242337, `RNS_PRIME_BITS'd501280585, `RNS_PRIME_BITS'd726033385, `RNS_PRIME_BITS'd915813205, `RNS_PRIME_BITS'd1232024916},
    '{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd755984682, `RNS_PRIME_BITS'd825850527, `RNS_PRIME_BITS'd867645482, `RNS_PRIME_BITS'd741438072, `RNS_PRIME_BITS'd1015419087, `RNS_PRIME_BITS'd1868974263, `RNS_PRIME_BITS'd1280052164, `RNS_PRIME_BITS'd576935286, `RNS_PRIME_BITS'd1803245003, `RNS_PRIME_BITS'd862452203},
    '{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd195958569, `RNS_PRIME_BITS'd1678176312, `RNS_PRIME_BITS'd1768673731, `RNS_PRIME_BITS'd377441427, `RNS_PRIME_BITS'd283910163, `RNS_PRIME_BITS'd714687244, `RNS_PRIME_BITS'd1414491618, `RNS_PRIME_BITS'd1114772995, `RNS_PRIME_BITS'd2038631761, `RNS_PRIME_BITS'd1235495758},
    '{`RNS_PRIME_BITS'd167, `RNS_PRIME_BITS'd711514739, `RNS_PRIME_BITS'd1837214212, `RNS_PRIME_BITS'd1945467504, `RNS_PRIME_BITS'd605421543, `RNS_PRIME_BITS'd558182534, `RNS_PRIME_BITS'd716094236, `RNS_PRIME_BITS'd1114379823, `RNS_PRIME_BITS'd271557768, `RNS_PRIME_BITS'd2097514289, `RNS_PRIME_BITS'd1782698780},
    '{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd707719628, `RNS_PRIME_BITS'd988967764, `RNS_PRIME_BITS'd2055368146, `RNS_PRIME_BITS'd1745192673, `RNS_PRIME_BITS'd177037800, `RNS_PRIME_BITS'd1835330505, `RNS_PRIME_BITS'd1017619763, `RNS_PRIME_BITS'd182878640, `RNS_PRIME_BITS'd546019738, `RNS_PRIME_BITS'd357572893}
};


const rns_residue_t A2__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1340328697, `RNS_PRIME_BITS'd1028411192, `RNS_PRIME_BITS'd833505390, `RNS_PRIME_BITS'd508914425, `RNS_PRIME_BITS'd695101177, `RNS_PRIME_BITS'd121929651, `RNS_PRIME_BITS'd468190141, `RNS_PRIME_BITS'd158621671, `RNS_PRIME_BITS'd1229496176, `RNS_PRIME_BITS'd1922507611},
    '{`RNS_PRIME_BITS'd227, `RNS_PRIME_BITS'd1897012015, `RNS_PRIME_BITS'd424664047, `RNS_PRIME_BITS'd148390489, `RNS_PRIME_BITS'd1660881012, `RNS_PRIME_BITS'd1839841661, `RNS_PRIME_BITS'd600890401, `RNS_PRIME_BITS'd111859334, `RNS_PRIME_BITS'd63012075, `RNS_PRIME_BITS'd1837715341, `RNS_PRIME_BITS'd2102711601},
    '{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd952024879, `RNS_PRIME_BITS'd1847294303, `RNS_PRIME_BITS'd1024507888, `RNS_PRIME_BITS'd1731714129, `RNS_PRIME_BITS'd456798983, `RNS_PRIME_BITS'd398357807, `RNS_PRIME_BITS'd819150038, `RNS_PRIME_BITS'd1074871179, `RNS_PRIME_BITS'd1881538838, `RNS_PRIME_BITS'd984786775},
    '{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd214890831, `RNS_PRIME_BITS'd1793609357, `RNS_PRIME_BITS'd293158148, `RNS_PRIME_BITS'd941952042, `RNS_PRIME_BITS'd1703338787, `RNS_PRIME_BITS'd477362987, `RNS_PRIME_BITS'd755957961, `RNS_PRIME_BITS'd1779634707, `RNS_PRIME_BITS'd886758664, `RNS_PRIME_BITS'd322190161},
    '{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd2013309932, `RNS_PRIME_BITS'd1196272423, `RNS_PRIME_BITS'd1913281042, `RNS_PRIME_BITS'd1933756359, `RNS_PRIME_BITS'd1005191015, `RNS_PRIME_BITS'd2100169185, `RNS_PRIME_BITS'd186901693, `RNS_PRIME_BITS'd1462544178, `RNS_PRIME_BITS'd642790623, `RNS_PRIME_BITS'd150495599},
    '{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd712620492, `RNS_PRIME_BITS'd253161811, `RNS_PRIME_BITS'd171550392, `RNS_PRIME_BITS'd2035805351, `RNS_PRIME_BITS'd2095024128, `RNS_PRIME_BITS'd1227883816, `RNS_PRIME_BITS'd575815669, `RNS_PRIME_BITS'd2002458832, `RNS_PRIME_BITS'd1563852721, `RNS_PRIME_BITS'd508758874},
    '{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd832585577, `RNS_PRIME_BITS'd357443542, `RNS_PRIME_BITS'd283467771, `RNS_PRIME_BITS'd856202594, `RNS_PRIME_BITS'd1002737735, `RNS_PRIME_BITS'd782790808, `RNS_PRIME_BITS'd1985333376, `RNS_PRIME_BITS'd245128879, `RNS_PRIME_BITS'd351791664, `RNS_PRIME_BITS'd1185501061},
    '{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd293386272, `RNS_PRIME_BITS'd1188507358, `RNS_PRIME_BITS'd22433621, `RNS_PRIME_BITS'd582320240, `RNS_PRIME_BITS'd2094628288, `RNS_PRIME_BITS'd828243241, `RNS_PRIME_BITS'd1318815447, `RNS_PRIME_BITS'd1561322294, `RNS_PRIME_BITS'd251856247, `RNS_PRIME_BITS'd586126026},
    '{`RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd707227732, `RNS_PRIME_BITS'd2074311491, `RNS_PRIME_BITS'd2131174023, `RNS_PRIME_BITS'd567084629, `RNS_PRIME_BITS'd1168712801, `RNS_PRIME_BITS'd1143862775, `RNS_PRIME_BITS'd399711304, `RNS_PRIME_BITS'd1164710298, `RNS_PRIME_BITS'd237095739, `RNS_PRIME_BITS'd1223221511},
    '{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd713648247, `RNS_PRIME_BITS'd479395508, `RNS_PRIME_BITS'd289517191, `RNS_PRIME_BITS'd270218379, `RNS_PRIME_BITS'd2100172118, `RNS_PRIME_BITS'd1611389917, `RNS_PRIME_BITS'd1301115129, `RNS_PRIME_BITS'd728629924, `RNS_PRIME_BITS'd1579218442, `RNS_PRIME_BITS'd271989711},
    '{`RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd237400224, `RNS_PRIME_BITS'd1139042970, `RNS_PRIME_BITS'd282688036, `RNS_PRIME_BITS'd869650008, `RNS_PRIME_BITS'd491537767, `RNS_PRIME_BITS'd1441081581, `RNS_PRIME_BITS'd655100268, `RNS_PRIME_BITS'd1557975835, `RNS_PRIME_BITS'd1026539034, `RNS_PRIME_BITS'd499527145},
    '{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd557753617, `RNS_PRIME_BITS'd878833429, `RNS_PRIME_BITS'd1373561798, `RNS_PRIME_BITS'd1844073307, `RNS_PRIME_BITS'd94445269, `RNS_PRIME_BITS'd2014326158, `RNS_PRIME_BITS'd343865196, `RNS_PRIME_BITS'd775191453, `RNS_PRIME_BITS'd1608547572, `RNS_PRIME_BITS'd126311803},
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd252932985, `RNS_PRIME_BITS'd1123198115, `RNS_PRIME_BITS'd896914588, `RNS_PRIME_BITS'd969680251, `RNS_PRIME_BITS'd1168800444, `RNS_PRIME_BITS'd1914069947, `RNS_PRIME_BITS'd263023560, `RNS_PRIME_BITS'd799316948, `RNS_PRIME_BITS'd352769466, `RNS_PRIME_BITS'd313895061},
    '{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd1771618026, `RNS_PRIME_BITS'd1407987179, `RNS_PRIME_BITS'd1723691945, `RNS_PRIME_BITS'd721970711, `RNS_PRIME_BITS'd1012620522, `RNS_PRIME_BITS'd404576311, `RNS_PRIME_BITS'd57230767, `RNS_PRIME_BITS'd1868541068, `RNS_PRIME_BITS'd1152816320, `RNS_PRIME_BITS'd621194939},
    '{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1242370691, `RNS_PRIME_BITS'd1436402501, `RNS_PRIME_BITS'd1305837762, `RNS_PRIME_BITS'd1420137746, `RNS_PRIME_BITS'd57070319, `RNS_PRIME_BITS'd1789467850, `RNS_PRIME_BITS'd586454966, `RNS_PRIME_BITS'd549398473, `RNS_PRIME_BITS'd595211950, `RNS_PRIME_BITS'd74535715},
    '{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd363925171, `RNS_PRIME_BITS'd1086348616, `RNS_PRIME_BITS'd353727616, `RNS_PRIME_BITS'd373279121, `RNS_PRIME_BITS'd518645799, `RNS_PRIME_BITS'd1473668681, `RNS_PRIME_BITS'd744013713, `RNS_PRIME_BITS'd629613559, `RNS_PRIME_BITS'd1943859100, `RNS_PRIME_BITS'd789731493},
    '{`RNS_PRIME_BITS'd230, `RNS_PRIME_BITS'd1218992033, `RNS_PRIME_BITS'd2056101164, `RNS_PRIME_BITS'd483236890, `RNS_PRIME_BITS'd347881410, `RNS_PRIME_BITS'd718379194, `RNS_PRIME_BITS'd89425199, `RNS_PRIME_BITS'd1226296273, `RNS_PRIME_BITS'd721891169, `RNS_PRIME_BITS'd2066476512, `RNS_PRIME_BITS'd1804991562},
    '{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd455237887, `RNS_PRIME_BITS'd1892988214, `RNS_PRIME_BITS'd1279868935, `RNS_PRIME_BITS'd603784556, `RNS_PRIME_BITS'd212834038, `RNS_PRIME_BITS'd492818166, `RNS_PRIME_BITS'd349005833, `RNS_PRIME_BITS'd856605567, `RNS_PRIME_BITS'd566636026, `RNS_PRIME_BITS'd200972298},
    '{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd352156915, `RNS_PRIME_BITS'd416537380, `RNS_PRIME_BITS'd2057979471, `RNS_PRIME_BITS'd521394630, `RNS_PRIME_BITS'd520005871, `RNS_PRIME_BITS'd1371324822, `RNS_PRIME_BITS'd95777377, `RNS_PRIME_BITS'd138940384, `RNS_PRIME_BITS'd1847750006, `RNS_PRIME_BITS'd626091291},
    '{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd1765902167, `RNS_PRIME_BITS'd237580393, `RNS_PRIME_BITS'd1583354238, `RNS_PRIME_BITS'd881356348, `RNS_PRIME_BITS'd55580668, `RNS_PRIME_BITS'd447871555, `RNS_PRIME_BITS'd495777285, `RNS_PRIME_BITS'd1402912932, `RNS_PRIME_BITS'd1589862690, `RNS_PRIME_BITS'd1961501413},
    '{`RNS_PRIME_BITS'd174, `RNS_PRIME_BITS'd452946413, `RNS_PRIME_BITS'd1648354070, `RNS_PRIME_BITS'd1953678431, `RNS_PRIME_BITS'd1895756983, `RNS_PRIME_BITS'd327607571, `RNS_PRIME_BITS'd306136394, `RNS_PRIME_BITS'd893032770, `RNS_PRIME_BITS'd1339902012, `RNS_PRIME_BITS'd907888793, `RNS_PRIME_BITS'd2096271269},
    '{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd530928021, `RNS_PRIME_BITS'd1045149885, `RNS_PRIME_BITS'd620184326, `RNS_PRIME_BITS'd1854123236, `RNS_PRIME_BITS'd164062551, `RNS_PRIME_BITS'd1709464154, `RNS_PRIME_BITS'd168182394, `RNS_PRIME_BITS'd334728737, `RNS_PRIME_BITS'd213279582, `RNS_PRIME_BITS'd1255432417},
    '{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd1202546534, `RNS_PRIME_BITS'd1254129065, `RNS_PRIME_BITS'd1579796147, `RNS_PRIME_BITS'd1787262223, `RNS_PRIME_BITS'd1705922028, `RNS_PRIME_BITS'd508253148, `RNS_PRIME_BITS'd1313033174, `RNS_PRIME_BITS'd807185662, `RNS_PRIME_BITS'd259916130, `RNS_PRIME_BITS'd456307767},
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd34800640, `RNS_PRIME_BITS'd1761558539, `RNS_PRIME_BITS'd228331537, `RNS_PRIME_BITS'd1422312480, `RNS_PRIME_BITS'd432608989, `RNS_PRIME_BITS'd1148635437, `RNS_PRIME_BITS'd1685559959, `RNS_PRIME_BITS'd1710561155, `RNS_PRIME_BITS'd670637027, `RNS_PRIME_BITS'd101903952},
    '{`RNS_PRIME_BITS'd38, `RNS_PRIME_BITS'd1563853717, `RNS_PRIME_BITS'd571201328, `RNS_PRIME_BITS'd245251714, `RNS_PRIME_BITS'd1663970889, `RNS_PRIME_BITS'd1902173506, `RNS_PRIME_BITS'd189846866, `RNS_PRIME_BITS'd1451639541, `RNS_PRIME_BITS'd1558590312, `RNS_PRIME_BITS'd2006475795, `RNS_PRIME_BITS'd731899446},
    '{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd953006543, `RNS_PRIME_BITS'd1333419366, `RNS_PRIME_BITS'd803996697, `RNS_PRIME_BITS'd699638571, `RNS_PRIME_BITS'd1570575928, `RNS_PRIME_BITS'd1754980088, `RNS_PRIME_BITS'd706796035, `RNS_PRIME_BITS'd1027625782, `RNS_PRIME_BITS'd2133888631, `RNS_PRIME_BITS'd1162595841},
    '{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd1637537897, `RNS_PRIME_BITS'd20482474, `RNS_PRIME_BITS'd889619225, `RNS_PRIME_BITS'd1780328347, `RNS_PRIME_BITS'd1517088642, `RNS_PRIME_BITS'd1435596795, `RNS_PRIME_BITS'd1930430867, `RNS_PRIME_BITS'd1520097171, `RNS_PRIME_BITS'd1029411705, `RNS_PRIME_BITS'd506584303},
    '{`RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd1518024326, `RNS_PRIME_BITS'd1927616150, `RNS_PRIME_BITS'd1161933470, `RNS_PRIME_BITS'd1072463355, `RNS_PRIME_BITS'd2079805121, `RNS_PRIME_BITS'd1570064471, `RNS_PRIME_BITS'd149929679, `RNS_PRIME_BITS'd306716022, `RNS_PRIME_BITS'd1496495185, `RNS_PRIME_BITS'd1041866057},
    '{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd1400343730, `RNS_PRIME_BITS'd32890735, `RNS_PRIME_BITS'd1645109039, `RNS_PRIME_BITS'd332720266, `RNS_PRIME_BITS'd522951379, `RNS_PRIME_BITS'd1266211659, `RNS_PRIME_BITS'd1374693309, `RNS_PRIME_BITS'd874681560, `RNS_PRIME_BITS'd204708434, `RNS_PRIME_BITS'd609873395},
    '{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd2117964355, `RNS_PRIME_BITS'd1542791771, `RNS_PRIME_BITS'd259735212, `RNS_PRIME_BITS'd1640745609, `RNS_PRIME_BITS'd1283940151, `RNS_PRIME_BITS'd929408010, `RNS_PRIME_BITS'd1005391845, `RNS_PRIME_BITS'd295962104, `RNS_PRIME_BITS'd18063076, `RNS_PRIME_BITS'd2128075980},
    '{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd1385643703, `RNS_PRIME_BITS'd726954292, `RNS_PRIME_BITS'd1736206351, `RNS_PRIME_BITS'd680972654, `RNS_PRIME_BITS'd1491864843, `RNS_PRIME_BITS'd930967383, `RNS_PRIME_BITS'd1412993692, `RNS_PRIME_BITS'd1701231324, `RNS_PRIME_BITS'd983954389, `RNS_PRIME_BITS'd775122167},
    '{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd682683785, `RNS_PRIME_BITS'd1458002286, `RNS_PRIME_BITS'd130064439, `RNS_PRIME_BITS'd515229608, `RNS_PRIME_BITS'd240014085, `RNS_PRIME_BITS'd732547739, `RNS_PRIME_BITS'd700413047, `RNS_PRIME_BITS'd1405345957, `RNS_PRIME_BITS'd290637115, `RNS_PRIME_BITS'd990713641},
    '{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd364431565, `RNS_PRIME_BITS'd1277017596, `RNS_PRIME_BITS'd1522582382, `RNS_PRIME_BITS'd1786416419, `RNS_PRIME_BITS'd861608707, `RNS_PRIME_BITS'd1284337464, `RNS_PRIME_BITS'd1071267324, `RNS_PRIME_BITS'd1115579539, `RNS_PRIME_BITS'd1943030248, `RNS_PRIME_BITS'd1035515045},
    '{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd1564900277, `RNS_PRIME_BITS'd672953399, `RNS_PRIME_BITS'd533116035, `RNS_PRIME_BITS'd1971824569, `RNS_PRIME_BITS'd256140759, `RNS_PRIME_BITS'd550284574, `RNS_PRIME_BITS'd1868169509, `RNS_PRIME_BITS'd1949422640, `RNS_PRIME_BITS'd787871302, `RNS_PRIME_BITS'd1915179667},
    '{`RNS_PRIME_BITS'd37, `RNS_PRIME_BITS'd888635231, `RNS_PRIME_BITS'd591286787, `RNS_PRIME_BITS'd2142481268, `RNS_PRIME_BITS'd2049260352, `RNS_PRIME_BITS'd1140808319, `RNS_PRIME_BITS'd321165315, `RNS_PRIME_BITS'd965976563, `RNS_PRIME_BITS'd1671350840, `RNS_PRIME_BITS'd1644418855, `RNS_PRIME_BITS'd1677324236},
    '{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd1637530535, `RNS_PRIME_BITS'd2087681052, `RNS_PRIME_BITS'd1478245845, `RNS_PRIME_BITS'd995137290, `RNS_PRIME_BITS'd584188626, `RNS_PRIME_BITS'd1885333088, `RNS_PRIME_BITS'd1845090887, `RNS_PRIME_BITS'd428160732, `RNS_PRIME_BITS'd1073719221, `RNS_PRIME_BITS'd1448512584},
    '{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd1749950010, `RNS_PRIME_BITS'd580420431, `RNS_PRIME_BITS'd892596393, `RNS_PRIME_BITS'd1019570997, `RNS_PRIME_BITS'd885458894, `RNS_PRIME_BITS'd514520152, `RNS_PRIME_BITS'd336938809, `RNS_PRIME_BITS'd1211993469, `RNS_PRIME_BITS'd630510729, `RNS_PRIME_BITS'd1561927548},
    '{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd387697373, `RNS_PRIME_BITS'd1513009803, `RNS_PRIME_BITS'd1122647403, `RNS_PRIME_BITS'd423356178, `RNS_PRIME_BITS'd732466220, `RNS_PRIME_BITS'd1449223682, `RNS_PRIME_BITS'd855139304, `RNS_PRIME_BITS'd1746389734, `RNS_PRIME_BITS'd1042485439, `RNS_PRIME_BITS'd965972923},
    '{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd1103034900, `RNS_PRIME_BITS'd187595593, `RNS_PRIME_BITS'd708552635, `RNS_PRIME_BITS'd195619786, `RNS_PRIME_BITS'd1776899433, `RNS_PRIME_BITS'd1897397501, `RNS_PRIME_BITS'd1883876023, `RNS_PRIME_BITS'd909312593, `RNS_PRIME_BITS'd1828144020, `RNS_PRIME_BITS'd1271430307},
    '{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd972408796, `RNS_PRIME_BITS'd1667335346, `RNS_PRIME_BITS'd1348489626, `RNS_PRIME_BITS'd1422461612, `RNS_PRIME_BITS'd1880010760, `RNS_PRIME_BITS'd423612396, `RNS_PRIME_BITS'd507740764, `RNS_PRIME_BITS'd144120395, `RNS_PRIME_BITS'd1318962956, `RNS_PRIME_BITS'd619499839},
    '{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd948585442, `RNS_PRIME_BITS'd13763333, `RNS_PRIME_BITS'd685888583, `RNS_PRIME_BITS'd169247853, `RNS_PRIME_BITS'd239620760, `RNS_PRIME_BITS'd725391476, `RNS_PRIME_BITS'd276938486, `RNS_PRIME_BITS'd488687644, `RNS_PRIME_BITS'd139413933, `RNS_PRIME_BITS'd556100233},
    '{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd455635859, `RNS_PRIME_BITS'd2046527541, `RNS_PRIME_BITS'd688338515, `RNS_PRIME_BITS'd789628807, `RNS_PRIME_BITS'd776121815, `RNS_PRIME_BITS'd2015930360, `RNS_PRIME_BITS'd1039112052, `RNS_PRIME_BITS'd1257796053, `RNS_PRIME_BITS'd1363141974, `RNS_PRIME_BITS'd1849975529},
    '{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1451617879, `RNS_PRIME_BITS'd911347881, `RNS_PRIME_BITS'd830018904, `RNS_PRIME_BITS'd1194628656, `RNS_PRIME_BITS'd1301376534, `RNS_PRIME_BITS'd2101833799, `RNS_PRIME_BITS'd1029298036, `RNS_PRIME_BITS'd934458470, `RNS_PRIME_BITS'd1434806506, `RNS_PRIME_BITS'd50832969},
    '{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1923221321, `RNS_PRIME_BITS'd574863860, `RNS_PRIME_BITS'd1825964470, `RNS_PRIME_BITS'd1080821454, `RNS_PRIME_BITS'd1628149686, `RNS_PRIME_BITS'd1111625142, `RNS_PRIME_BITS'd1967290119, `RNS_PRIME_BITS'd963652876, `RNS_PRIME_BITS'd693488822, `RNS_PRIME_BITS'd936107445},
    '{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd1239035345, `RNS_PRIME_BITS'd1396123321, `RNS_PRIME_BITS'd649161926, `RNS_PRIME_BITS'd597549788, `RNS_PRIME_BITS'd807581434, `RNS_PRIME_BITS'd1657302521, `RNS_PRIME_BITS'd350202451, `RNS_PRIME_BITS'd1469810176, `RNS_PRIME_BITS'd1731537838, `RNS_PRIME_BITS'd1473677131},
    '{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd1927225614, `RNS_PRIME_BITS'd169557685, `RNS_PRIME_BITS'd1124531029, `RNS_PRIME_BITS'd645893142, `RNS_PRIME_BITS'd11808009, `RNS_PRIME_BITS'd1318488075, `RNS_PRIME_BITS'd399784272, `RNS_PRIME_BITS'd935117004, `RNS_PRIME_BITS'd787168005, `RNS_PRIME_BITS'd1311169409},
    '{`RNS_PRIME_BITS'd179, `RNS_PRIME_BITS'd854068432, `RNS_PRIME_BITS'd320347225, `RNS_PRIME_BITS'd1658503202, `RNS_PRIME_BITS'd127165862, `RNS_PRIME_BITS'd578927198, `RNS_PRIME_BITS'd766179215, `RNS_PRIME_BITS'd1048877454, `RNS_PRIME_BITS'd941095724, `RNS_PRIME_BITS'd956202953, `RNS_PRIME_BITS'd1293147664},
    '{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd678560121, `RNS_PRIME_BITS'd2109389178, `RNS_PRIME_BITS'd1643846849, `RNS_PRIME_BITS'd1393021507, `RNS_PRIME_BITS'd1923080752, `RNS_PRIME_BITS'd576549368, `RNS_PRIME_BITS'd1256355067, `RNS_PRIME_BITS'd950129201, `RNS_PRIME_BITS'd1498451417, `RNS_PRIME_BITS'd1529713522},
    '{`RNS_PRIME_BITS'd233, `RNS_PRIME_BITS'd485324390, `RNS_PRIME_BITS'd867109936, `RNS_PRIME_BITS'd614876355, `RNS_PRIME_BITS'd813104772, `RNS_PRIME_BITS'd2014655754, `RNS_PRIME_BITS'd579028278, `RNS_PRIME_BITS'd637212477, `RNS_PRIME_BITS'd1457836900, `RNS_PRIME_BITS'd936084674, `RNS_PRIME_BITS'd1257556765},
    '{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd1270140768, `RNS_PRIME_BITS'd289457166, `RNS_PRIME_BITS'd636248138, `RNS_PRIME_BITS'd420615460, `RNS_PRIME_BITS'd1080981210, `RNS_PRIME_BITS'd1715305531, `RNS_PRIME_BITS'd865940732, `RNS_PRIME_BITS'd1181573363, `RNS_PRIME_BITS'd85644503, `RNS_PRIME_BITS'd1563555965},
    '{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd605171683, `RNS_PRIME_BITS'd935946349, `RNS_PRIME_BITS'd934562408, `RNS_PRIME_BITS'd692311391, `RNS_PRIME_BITS'd2129468798, `RNS_PRIME_BITS'd492377783, `RNS_PRIME_BITS'd370107380, `RNS_PRIME_BITS'd1734485218, `RNS_PRIME_BITS'd1953235194, `RNS_PRIME_BITS'd12929148},
    '{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd845066254, `RNS_PRIME_BITS'd383929236, `RNS_PRIME_BITS'd1727537090, `RNS_PRIME_BITS'd524673580, `RNS_PRIME_BITS'd1110222294, `RNS_PRIME_BITS'd942316711, `RNS_PRIME_BITS'd710838697, `RNS_PRIME_BITS'd881641935, `RNS_PRIME_BITS'd1476192243, `RNS_PRIME_BITS'd1301340958},
    '{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd523124056, `RNS_PRIME_BITS'd1725990315, `RNS_PRIME_BITS'd1802356227, `RNS_PRIME_BITS'd929179022, `RNS_PRIME_BITS'd2038391289, `RNS_PRIME_BITS'd763417140, `RNS_PRIME_BITS'd1867905882, `RNS_PRIME_BITS'd240396442, `RNS_PRIME_BITS'd1514687753, `RNS_PRIME_BITS'd662086514},
    '{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd1008923926, `RNS_PRIME_BITS'd1712267184, `RNS_PRIME_BITS'd66715980, `RNS_PRIME_BITS'd2116786604, `RNS_PRIME_BITS'd1705268748, `RNS_PRIME_BITS'd167592567, `RNS_PRIME_BITS'd941595340, `RNS_PRIME_BITS'd2112950272, `RNS_PRIME_BITS'd966183466, `RNS_PRIME_BITS'd68405799},
    '{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd303034312, `RNS_PRIME_BITS'd125642853, `RNS_PRIME_BITS'd1409626079, `RNS_PRIME_BITS'd1641311794, `RNS_PRIME_BITS'd943835740, `RNS_PRIME_BITS'd1569241352, `RNS_PRIME_BITS'd742445703, `RNS_PRIME_BITS'd1396267602, `RNS_PRIME_BITS'd62563416, `RNS_PRIME_BITS'd359370362},
    '{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd1751464864, `RNS_PRIME_BITS'd523326004, `RNS_PRIME_BITS'd1335530113, `RNS_PRIME_BITS'd765454914, `RNS_PRIME_BITS'd1668622198, `RNS_PRIME_BITS'd117421188, `RNS_PRIME_BITS'd1924208047, `RNS_PRIME_BITS'd1595402938, `RNS_PRIME_BITS'd1870251196, `RNS_PRIME_BITS'd1067446201},
    '{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd1580803029, `RNS_PRIME_BITS'd176956725, `RNS_PRIME_BITS'd1091609407, `RNS_PRIME_BITS'd1945581937, `RNS_PRIME_BITS'd1758300001, `RNS_PRIME_BITS'd350292717, `RNS_PRIME_BITS'd1114617248, `RNS_PRIME_BITS'd590064287, `RNS_PRIME_BITS'd986480542, `RNS_PRIME_BITS'd424378780},
    '{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd97191010, `RNS_PRIME_BITS'd1363669740, `RNS_PRIME_BITS'd668503916, `RNS_PRIME_BITS'd500864865, `RNS_PRIME_BITS'd631297502, `RNS_PRIME_BITS'd1109658718, `RNS_PRIME_BITS'd532533810, `RNS_PRIME_BITS'd936353871, `RNS_PRIME_BITS'd936998295, `RNS_PRIME_BITS'd2130785219},
    '{`RNS_PRIME_BITS'd151, `RNS_PRIME_BITS'd816211149, `RNS_PRIME_BITS'd1584074260, `RNS_PRIME_BITS'd1752514649, `RNS_PRIME_BITS'd1081668837, `RNS_PRIME_BITS'd474083483, `RNS_PRIME_BITS'd1356426305, `RNS_PRIME_BITS'd1086476956, `RNS_PRIME_BITS'd1019470604, `RNS_PRIME_BITS'd1037006672, `RNS_PRIME_BITS'd861969653},
    '{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1595186567, `RNS_PRIME_BITS'd1432874892, `RNS_PRIME_BITS'd1786110961, `RNS_PRIME_BITS'd1106254626, `RNS_PRIME_BITS'd1259076666, `RNS_PRIME_BITS'd1345402623, `RNS_PRIME_BITS'd119932553, `RNS_PRIME_BITS'd1067721364, `RNS_PRIME_BITS'd1368327433, `RNS_PRIME_BITS'd2145273054},
    '{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd1881822655, `RNS_PRIME_BITS'd1087427362, `RNS_PRIME_BITS'd1453347102, `RNS_PRIME_BITS'd1629269185, `RNS_PRIME_BITS'd1625128790, `RNS_PRIME_BITS'd1399142330, `RNS_PRIME_BITS'd124806697, `RNS_PRIME_BITS'd2128518943, `RNS_PRIME_BITS'd835731850, `RNS_PRIME_BITS'd1040493708},
    '{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd404944566, `RNS_PRIME_BITS'd329289509, `RNS_PRIME_BITS'd1147166527, `RNS_PRIME_BITS'd1500208368, `RNS_PRIME_BITS'd1075924044, `RNS_PRIME_BITS'd818763913, `RNS_PRIME_BITS'd2041605630, `RNS_PRIME_BITS'd33458838, `RNS_PRIME_BITS'd1105837464, `RNS_PRIME_BITS'd1741403262},
    '{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd466007139, `RNS_PRIME_BITS'd2085642063, `RNS_PRIME_BITS'd902279933, `RNS_PRIME_BITS'd930674557, `RNS_PRIME_BITS'd843689752, `RNS_PRIME_BITS'd723893333, `RNS_PRIME_BITS'd293672503, `RNS_PRIME_BITS'd1732507925, `RNS_PRIME_BITS'd1973944467, `RNS_PRIME_BITS'd298255786},
    '{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd1459654781, `RNS_PRIME_BITS'd914457688, `RNS_PRIME_BITS'd1441067476, `RNS_PRIME_BITS'd623050342, `RNS_PRIME_BITS'd1556747181, `RNS_PRIME_BITS'd1135592291, `RNS_PRIME_BITS'd1024092932, `RNS_PRIME_BITS'd998978140, `RNS_PRIME_BITS'd652166025, `RNS_PRIME_BITS'd1674169521}
};


const rns_residue_t B2__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd819594541, `RNS_PRIME_BITS'd634162875, `RNS_PRIME_BITS'd416060616, `RNS_PRIME_BITS'd1154266234, `RNS_PRIME_BITS'd264646753, `RNS_PRIME_BITS'd1294044377, `RNS_PRIME_BITS'd950158574, `RNS_PRIME_BITS'd1513440422, `RNS_PRIME_BITS'd510797271, `RNS_PRIME_BITS'd489440472},
    '{`RNS_PRIME_BITS'd201, `RNS_PRIME_BITS'd2099677320, `RNS_PRIME_BITS'd1394874675, `RNS_PRIME_BITS'd246679523, `RNS_PRIME_BITS'd147367499, `RNS_PRIME_BITS'd1043590720, `RNS_PRIME_BITS'd1582511291, `RNS_PRIME_BITS'd1209090269, `RNS_PRIME_BITS'd612566604, `RNS_PRIME_BITS'd738619560, `RNS_PRIME_BITS'd1179291959},
    '{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd258927414, `RNS_PRIME_BITS'd1564853585, `RNS_PRIME_BITS'd2019452836, `RNS_PRIME_BITS'd891764882, `RNS_PRIME_BITS'd1359612793, `RNS_PRIME_BITS'd1482587555, `RNS_PRIME_BITS'd797572148, `RNS_PRIME_BITS'd477094658, `RNS_PRIME_BITS'd326608941, `RNS_PRIME_BITS'd640982480},
    '{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd739401345, `RNS_PRIME_BITS'd1929523713, `RNS_PRIME_BITS'd1400841295, `RNS_PRIME_BITS'd770807619, `RNS_PRIME_BITS'd462147962, `RNS_PRIME_BITS'd1562561273, `RNS_PRIME_BITS'd1205264552, `RNS_PRIME_BITS'd1044595844, `RNS_PRIME_BITS'd1251653043, `RNS_PRIME_BITS'd552842898},
    '{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd1247659774, `RNS_PRIME_BITS'd391309228, `RNS_PRIME_BITS'd1024538162, `RNS_PRIME_BITS'd1791655406, `RNS_PRIME_BITS'd2080402555, `RNS_PRIME_BITS'd1666855140, `RNS_PRIME_BITS'd1927242802, `RNS_PRIME_BITS'd1064001599, `RNS_PRIME_BITS'd1912116412, `RNS_PRIME_BITS'd1169633428},
    '{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd1911121267, `RNS_PRIME_BITS'd705622761, `RNS_PRIME_BITS'd739670039, `RNS_PRIME_BITS'd909302999, `RNS_PRIME_BITS'd148429630, `RNS_PRIME_BITS'd826775931, `RNS_PRIME_BITS'd799157590, `RNS_PRIME_BITS'd878768208, `RNS_PRIME_BITS'd1549848748, `RNS_PRIME_BITS'd1203674672},
    '{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd2063930117, `RNS_PRIME_BITS'd1239914682, `RNS_PRIME_BITS'd1512585478, `RNS_PRIME_BITS'd767597841, `RNS_PRIME_BITS'd14632488, `RNS_PRIME_BITS'd944296056, `RNS_PRIME_BITS'd794245831, `RNS_PRIME_BITS'd1818032963, `RNS_PRIME_BITS'd865915820, `RNS_PRIME_BITS'd1353149695},
    '{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd2137032594, `RNS_PRIME_BITS'd160694812, `RNS_PRIME_BITS'd2042135464, `RNS_PRIME_BITS'd96815554, `RNS_PRIME_BITS'd1708371854, `RNS_PRIME_BITS'd2064372186, `RNS_PRIME_BITS'd231545040, `RNS_PRIME_BITS'd802166272, `RNS_PRIME_BITS'd1163026015, `RNS_PRIME_BITS'd1492809668},
    '{`RNS_PRIME_BITS'd167, `RNS_PRIME_BITS'd585108950, `RNS_PRIME_BITS'd1637316132, `RNS_PRIME_BITS'd1939982993, `RNS_PRIME_BITS'd551816934, `RNS_PRIME_BITS'd601710523, `RNS_PRIME_BITS'd500571176, `RNS_PRIME_BITS'd1262582881, `RNS_PRIME_BITS'd2128675054, `RNS_PRIME_BITS'd1432919089, `RNS_PRIME_BITS'd71493684},
    '{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd915546310, `RNS_PRIME_BITS'd1769984114, `RNS_PRIME_BITS'd1634450515, `RNS_PRIME_BITS'd1592951774, `RNS_PRIME_BITS'd1705215503, `RNS_PRIME_BITS'd1810505393, `RNS_PRIME_BITS'd344265867, `RNS_PRIME_BITS'd362893883, `RNS_PRIME_BITS'd773437356, `RNS_PRIME_BITS'd1541030357},
    '{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd320023023, `RNS_PRIME_BITS'd1633694795, `RNS_PRIME_BITS'd1277232447, `RNS_PRIME_BITS'd1214945910, `RNS_PRIME_BITS'd1290607431, `RNS_PRIME_BITS'd369284064, `RNS_PRIME_BITS'd1622292501, `RNS_PRIME_BITS'd590955314, `RNS_PRIME_BITS'd342395328, `RNS_PRIME_BITS'd685387560},
    '{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd63805057, `RNS_PRIME_BITS'd162020279, `RNS_PRIME_BITS'd1079972614, `RNS_PRIME_BITS'd1074912742, `RNS_PRIME_BITS'd320186892, `RNS_PRIME_BITS'd1081964391, `RNS_PRIME_BITS'd306135783, `RNS_PRIME_BITS'd748725398, `RNS_PRIME_BITS'd1357489485, `RNS_PRIME_BITS'd27601784},
    '{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd915789618, `RNS_PRIME_BITS'd492156747, `RNS_PRIME_BITS'd1890560517, `RNS_PRIME_BITS'd1499642241, `RNS_PRIME_BITS'd738472916, `RNS_PRIME_BITS'd1217845944, `RNS_PRIME_BITS'd9513635, `RNS_PRIME_BITS'd302480997, `RNS_PRIME_BITS'd429401349, `RNS_PRIME_BITS'd791717473},
    '{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd900496018, `RNS_PRIME_BITS'd1821279817, `RNS_PRIME_BITS'd370179856, `RNS_PRIME_BITS'd2091846937, `RNS_PRIME_BITS'd1733497094, `RNS_PRIME_BITS'd1454806983, `RNS_PRIME_BITS'd1911927544, `RNS_PRIME_BITS'd123883021, `RNS_PRIME_BITS'd403362422, `RNS_PRIME_BITS'd516266980},
    '{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd187169408, `RNS_PRIME_BITS'd527880281, `RNS_PRIME_BITS'd1404867017, `RNS_PRIME_BITS'd2094678075, `RNS_PRIME_BITS'd235416160, `RNS_PRIME_BITS'd1268826050, `RNS_PRIME_BITS'd750702119, `RNS_PRIME_BITS'd1107019521, `RNS_PRIME_BITS'd1188608593, `RNS_PRIME_BITS'd1424694820},
    '{`RNS_PRIME_BITS'd163, `RNS_PRIME_BITS'd1962284188, `RNS_PRIME_BITS'd405995600, `RNS_PRIME_BITS'd1860144132, `RNS_PRIME_BITS'd798327846, `RNS_PRIME_BITS'd1226026096, `RNS_PRIME_BITS'd183579250, `RNS_PRIME_BITS'd371890940, `RNS_PRIME_BITS'd1273651217, `RNS_PRIME_BITS'd1507770631, `RNS_PRIME_BITS'd1014435353},
    '{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd434472083, `RNS_PRIME_BITS'd1195837800, `RNS_PRIME_BITS'd2103407449, `RNS_PRIME_BITS'd1965061855, `RNS_PRIME_BITS'd206649400, `RNS_PRIME_BITS'd847617629, `RNS_PRIME_BITS'd542249444, `RNS_PRIME_BITS'd398466813, `RNS_PRIME_BITS'd452142554, `RNS_PRIME_BITS'd1994865915},
    '{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1708886127, `RNS_PRIME_BITS'd21734106, `RNS_PRIME_BITS'd1644786709, `RNS_PRIME_BITS'd1133762072, `RNS_PRIME_BITS'd101403870, `RNS_PRIME_BITS'd626538052, `RNS_PRIME_BITS'd63595079, `RNS_PRIME_BITS'd401308504, `RNS_PRIME_BITS'd708118132, `RNS_PRIME_BITS'd1141714988},
    '{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1406336163, `RNS_PRIME_BITS'd917044915, `RNS_PRIME_BITS'd1784945458, `RNS_PRIME_BITS'd1807509622, `RNS_PRIME_BITS'd1618340064, `RNS_PRIME_BITS'd2056570318, `RNS_PRIME_BITS'd1257821790, `RNS_PRIME_BITS'd125273275, `RNS_PRIME_BITS'd940657878, `RNS_PRIME_BITS'd370317992},
    '{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd2114345676, `RNS_PRIME_BITS'd755890229, `RNS_PRIME_BITS'd1785417238, `RNS_PRIME_BITS'd433814653, `RNS_PRIME_BITS'd1826163058, `RNS_PRIME_BITS'd1211851382, `RNS_PRIME_BITS'd432931088, `RNS_PRIME_BITS'd2102654617, `RNS_PRIME_BITS'd1337902533, `RNS_PRIME_BITS'd1923230210},
    '{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd1764916303, `RNS_PRIME_BITS'd204792833, `RNS_PRIME_BITS'd1529220788, `RNS_PRIME_BITS'd754892119, `RNS_PRIME_BITS'd1233638850, `RNS_PRIME_BITS'd539059468, `RNS_PRIME_BITS'd950427989, `RNS_PRIME_BITS'd1300131393, `RNS_PRIME_BITS'd1911425272, `RNS_PRIME_BITS'd1046872351},
    '{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd795705422, `RNS_PRIME_BITS'd307112129, `RNS_PRIME_BITS'd578197630, `RNS_PRIME_BITS'd790226394, `RNS_PRIME_BITS'd686008000, `RNS_PRIME_BITS'd310783029, `RNS_PRIME_BITS'd2105070156, `RNS_PRIME_BITS'd61914444, `RNS_PRIME_BITS'd1530203265, `RNS_PRIME_BITS'd343976073},
    '{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd649620690, `RNS_PRIME_BITS'd290477271, `RNS_PRIME_BITS'd814298234, `RNS_PRIME_BITS'd797115477, `RNS_PRIME_BITS'd1141346910, `RNS_PRIME_BITS'd585449069, `RNS_PRIME_BITS'd1627518941, `RNS_PRIME_BITS'd207871774, `RNS_PRIME_BITS'd157538684, `RNS_PRIME_BITS'd589066519},
    '{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd10593591, `RNS_PRIME_BITS'd1315039663, `RNS_PRIME_BITS'd1711382794, `RNS_PRIME_BITS'd1379485415, `RNS_PRIME_BITS'd1640851746, `RNS_PRIME_BITS'd1136932273, `RNS_PRIME_BITS'd423568379, `RNS_PRIME_BITS'd773279288, `RNS_PRIME_BITS'd1580401593, `RNS_PRIME_BITS'd990756297},
    '{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd1037357647, `RNS_PRIME_BITS'd1880641985, `RNS_PRIME_BITS'd1815670141, `RNS_PRIME_BITS'd811775812, `RNS_PRIME_BITS'd383333173, `RNS_PRIME_BITS'd1925215314, `RNS_PRIME_BITS'd515541833, `RNS_PRIME_BITS'd911697722, `RNS_PRIME_BITS'd1950762573, `RNS_PRIME_BITS'd2106453894},
    '{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd505170994, `RNS_PRIME_BITS'd1989781486, `RNS_PRIME_BITS'd1856998027, `RNS_PRIME_BITS'd322222698, `RNS_PRIME_BITS'd1120433740, `RNS_PRIME_BITS'd906370741, `RNS_PRIME_BITS'd40538345, `RNS_PRIME_BITS'd1546724914, `RNS_PRIME_BITS'd440647084, `RNS_PRIME_BITS'd608733417},
    '{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd45183827, `RNS_PRIME_BITS'd1871540698, `RNS_PRIME_BITS'd2016433637, `RNS_PRIME_BITS'd1839729940, `RNS_PRIME_BITS'd1995915962, `RNS_PRIME_BITS'd359544319, `RNS_PRIME_BITS'd958241987, `RNS_PRIME_BITS'd1899818794, `RNS_PRIME_BITS'd1389431075, `RNS_PRIME_BITS'd514254217},
    '{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd808516533, `RNS_PRIME_BITS'd288108504, `RNS_PRIME_BITS'd1779630901, `RNS_PRIME_BITS'd251205848, `RNS_PRIME_BITS'd1332817228, `RNS_PRIME_BITS'd871687548, `RNS_PRIME_BITS'd537877348, `RNS_PRIME_BITS'd1815713408, `RNS_PRIME_BITS'd1927809612, `RNS_PRIME_BITS'd2002278687},
    '{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd1683576530, `RNS_PRIME_BITS'd691310118, `RNS_PRIME_BITS'd9759421, `RNS_PRIME_BITS'd315304674, `RNS_PRIME_BITS'd1501326164, `RNS_PRIME_BITS'd1343653819, `RNS_PRIME_BITS'd62806841, `RNS_PRIME_BITS'd1479987306, `RNS_PRIME_BITS'd408322850, `RNS_PRIME_BITS'd15854668},
    '{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd685522807, `RNS_PRIME_BITS'd1850961964, `RNS_PRIME_BITS'd1338318113, `RNS_PRIME_BITS'd1173062040, `RNS_PRIME_BITS'd926763893, `RNS_PRIME_BITS'd219410216, `RNS_PRIME_BITS'd487931557, `RNS_PRIME_BITS'd682918185, `RNS_PRIME_BITS'd230619592, `RNS_PRIME_BITS'd1000310103},
    '{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1167225490, `RNS_PRIME_BITS'd525385688, `RNS_PRIME_BITS'd1745161141, `RNS_PRIME_BITS'd2092847354, `RNS_PRIME_BITS'd892798744, `RNS_PRIME_BITS'd1401580004, `RNS_PRIME_BITS'd1011219402, `RNS_PRIME_BITS'd465573817, `RNS_PRIME_BITS'd129325776, `RNS_PRIME_BITS'd1071014226},
    '{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd507364864, `RNS_PRIME_BITS'd1563159290, `RNS_PRIME_BITS'd1365781817, `RNS_PRIME_BITS'd63469545, `RNS_PRIME_BITS'd1075610931, `RNS_PRIME_BITS'd1984736416, `RNS_PRIME_BITS'd1421309240, `RNS_PRIME_BITS'd908302735, `RNS_PRIME_BITS'd1952866777, `RNS_PRIME_BITS'd1659354015},
    '{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd1850216089, `RNS_PRIME_BITS'd1876205824, `RNS_PRIME_BITS'd1909699201, `RNS_PRIME_BITS'd232283773, `RNS_PRIME_BITS'd315223926, `RNS_PRIME_BITS'd1778499474, `RNS_PRIME_BITS'd865164275, `RNS_PRIME_BITS'd1679998136, `RNS_PRIME_BITS'd759745972, `RNS_PRIME_BITS'd656494697},
    '{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1865733027, `RNS_PRIME_BITS'd667006867, `RNS_PRIME_BITS'd835234463, `RNS_PRIME_BITS'd2082753757, `RNS_PRIME_BITS'd760281410, `RNS_PRIME_BITS'd135500265, `RNS_PRIME_BITS'd1608769801, `RNS_PRIME_BITS'd514408626, `RNS_PRIME_BITS'd659313085, `RNS_PRIME_BITS'd1310779779},
    '{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1259530563, `RNS_PRIME_BITS'd476318156, `RNS_PRIME_BITS'd680762550, `RNS_PRIME_BITS'd159981766, `RNS_PRIME_BITS'd2033001506, `RNS_PRIME_BITS'd229622041, `RNS_PRIME_BITS'd509257478, `RNS_PRIME_BITS'd543362069, `RNS_PRIME_BITS'd103697047, `RNS_PRIME_BITS'd469819335},
    '{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd1937543422, `RNS_PRIME_BITS'd1584544453, `RNS_PRIME_BITS'd1030079444, `RNS_PRIME_BITS'd1581533698, `RNS_PRIME_BITS'd287727089, `RNS_PRIME_BITS'd1383795099, `RNS_PRIME_BITS'd1357499876, `RNS_PRIME_BITS'd2101530143, `RNS_PRIME_BITS'd2109492612, `RNS_PRIME_BITS'd344117895},
    '{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1588040718, `RNS_PRIME_BITS'd581138960, `RNS_PRIME_BITS'd374659106, `RNS_PRIME_BITS'd1499255422, `RNS_PRIME_BITS'd1646577730, `RNS_PRIME_BITS'd1573543715, `RNS_PRIME_BITS'd61131978, `RNS_PRIME_BITS'd1228581758, `RNS_PRIME_BITS'd635041661, `RNS_PRIME_BITS'd1074368433},
    '{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd353151117, `RNS_PRIME_BITS'd1901108366, `RNS_PRIME_BITS'd242482367, `RNS_PRIME_BITS'd519832032, `RNS_PRIME_BITS'd1392418783, `RNS_PRIME_BITS'd62306134, `RNS_PRIME_BITS'd1941131410, `RNS_PRIME_BITS'd1942740237, `RNS_PRIME_BITS'd563391763, `RNS_PRIME_BITS'd413079716},
    '{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd1512092102, `RNS_PRIME_BITS'd1004993657, `RNS_PRIME_BITS'd370115865, `RNS_PRIME_BITS'd1875428203, `RNS_PRIME_BITS'd1497052945, `RNS_PRIME_BITS'd1585766741, `RNS_PRIME_BITS'd1412955170, `RNS_PRIME_BITS'd501302283, `RNS_PRIME_BITS'd702748574, `RNS_PRIME_BITS'd1225237195},
    '{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd520149647, `RNS_PRIME_BITS'd515840591, `RNS_PRIME_BITS'd1498299651, `RNS_PRIME_BITS'd951545154, `RNS_PRIME_BITS'd639081141, `RNS_PRIME_BITS'd1059491839, `RNS_PRIME_BITS'd747090048, `RNS_PRIME_BITS'd1961143623, `RNS_PRIME_BITS'd400265686, `RNS_PRIME_BITS'd1198064782},
    '{`RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd1633012317, `RNS_PRIME_BITS'd1899398374, `RNS_PRIME_BITS'd128854806, `RNS_PRIME_BITS'd837024258, `RNS_PRIME_BITS'd2036820034, `RNS_PRIME_BITS'd1415002189, `RNS_PRIME_BITS'd553634427, `RNS_PRIME_BITS'd2076305601, `RNS_PRIME_BITS'd76323295, `RNS_PRIME_BITS'd414637077},
    '{`RNS_PRIME_BITS'd238, `RNS_PRIME_BITS'd1349680491, `RNS_PRIME_BITS'd1885788376, `RNS_PRIME_BITS'd2095417361, `RNS_PRIME_BITS'd1119908857, `RNS_PRIME_BITS'd1421065111, `RNS_PRIME_BITS'd1223027883, `RNS_PRIME_BITS'd151382370, `RNS_PRIME_BITS'd436880577, `RNS_PRIME_BITS'd1046791116, `RNS_PRIME_BITS'd1925704258},
    '{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1485058326, `RNS_PRIME_BITS'd163218604, `RNS_PRIME_BITS'd362222291, `RNS_PRIME_BITS'd2089249362, `RNS_PRIME_BITS'd1783759357, `RNS_PRIME_BITS'd467135732, `RNS_PRIME_BITS'd1902375748, `RNS_PRIME_BITS'd543808913, `RNS_PRIME_BITS'd248239272, `RNS_PRIME_BITS'd1626540682},
    '{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd2071347512, `RNS_PRIME_BITS'd1236608506, `RNS_PRIME_BITS'd1737180624, `RNS_PRIME_BITS'd1222965152, `RNS_PRIME_BITS'd1691308328, `RNS_PRIME_BITS'd1113227518, `RNS_PRIME_BITS'd2001857041, `RNS_PRIME_BITS'd1918939871, `RNS_PRIME_BITS'd860140296, `RNS_PRIME_BITS'd1495208452},
    '{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd1791435174, `RNS_PRIME_BITS'd1084854030, `RNS_PRIME_BITS'd621860874, `RNS_PRIME_BITS'd1847956270, `RNS_PRIME_BITS'd1433278422, `RNS_PRIME_BITS'd2015090342, `RNS_PRIME_BITS'd1140134113, `RNS_PRIME_BITS'd387546390, `RNS_PRIME_BITS'd1875855755, `RNS_PRIME_BITS'd1826620531},
    '{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd1969319885, `RNS_PRIME_BITS'd1216157117, `RNS_PRIME_BITS'd730992467, `RNS_PRIME_BITS'd1878086538, `RNS_PRIME_BITS'd1020341647, `RNS_PRIME_BITS'd499438714, `RNS_PRIME_BITS'd1809855918, `RNS_PRIME_BITS'd1385221753, `RNS_PRIME_BITS'd1961683318, `RNS_PRIME_BITS'd37117288},
    '{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd1239046013, `RNS_PRIME_BITS'd721545417, `RNS_PRIME_BITS'd884781361, `RNS_PRIME_BITS'd2141877786, `RNS_PRIME_BITS'd506316101, `RNS_PRIME_BITS'd470970922, `RNS_PRIME_BITS'd1225090919, `RNS_PRIME_BITS'd718658588, `RNS_PRIME_BITS'd1568470192, `RNS_PRIME_BITS'd1664245285},
    '{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd2073859149, `RNS_PRIME_BITS'd489244136, `RNS_PRIME_BITS'd559889519, `RNS_PRIME_BITS'd1182433981, `RNS_PRIME_BITS'd2031475892, `RNS_PRIME_BITS'd42550270, `RNS_PRIME_BITS'd1842190455, `RNS_PRIME_BITS'd807987319, `RNS_PRIME_BITS'd269870558, `RNS_PRIME_BITS'd271371964},
    '{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd984322734, `RNS_PRIME_BITS'd824282316, `RNS_PRIME_BITS'd112237508, `RNS_PRIME_BITS'd281203694, `RNS_PRIME_BITS'd1042679965, `RNS_PRIME_BITS'd534649879, `RNS_PRIME_BITS'd973730440, `RNS_PRIME_BITS'd587091442, `RNS_PRIME_BITS'd519490093, `RNS_PRIME_BITS'd35005606},
    '{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd1630999126, `RNS_PRIME_BITS'd340531089, `RNS_PRIME_BITS'd1688081553, `RNS_PRIME_BITS'd385333044, `RNS_PRIME_BITS'd1878325669, `RNS_PRIME_BITS'd1633392792, `RNS_PRIME_BITS'd1807393328, `RNS_PRIME_BITS'd595045519, `RNS_PRIME_BITS'd1613425123, `RNS_PRIME_BITS'd219343411},
    '{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd36729657, `RNS_PRIME_BITS'd1508989410, `RNS_PRIME_BITS'd1830400439, `RNS_PRIME_BITS'd82583994, `RNS_PRIME_BITS'd1805805965, `RNS_PRIME_BITS'd196658475, `RNS_PRIME_BITS'd278215989, `RNS_PRIME_BITS'd2138056788, `RNS_PRIME_BITS'd1724214718, `RNS_PRIME_BITS'd1600476637},
    '{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd918617112, `RNS_PRIME_BITS'd557513935, `RNS_PRIME_BITS'd937998310, `RNS_PRIME_BITS'd157008109, `RNS_PRIME_BITS'd1422187124, `RNS_PRIME_BITS'd1083468849, `RNS_PRIME_BITS'd1192876942, `RNS_PRIME_BITS'd1579861561, `RNS_PRIME_BITS'd311266371, `RNS_PRIME_BITS'd1598272211},
    '{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd1619949148, `RNS_PRIME_BITS'd1869077212, `RNS_PRIME_BITS'd1052858990, `RNS_PRIME_BITS'd1983164030, `RNS_PRIME_BITS'd460623130, `RNS_PRIME_BITS'd908142441, `RNS_PRIME_BITS'd435004017, `RNS_PRIME_BITS'd789128822, `RNS_PRIME_BITS'd623154567, `RNS_PRIME_BITS'd475302146},
    '{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd1254656805, `RNS_PRIME_BITS'd939423614, `RNS_PRIME_BITS'd217426264, `RNS_PRIME_BITS'd793662264, `RNS_PRIME_BITS'd1438970054, `RNS_PRIME_BITS'd1813246672, `RNS_PRIME_BITS'd1760659137, `RNS_PRIME_BITS'd1610565969, `RNS_PRIME_BITS'd669839356, `RNS_PRIME_BITS'd515008054},
    '{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd801292754, `RNS_PRIME_BITS'd125414131, `RNS_PRIME_BITS'd1835109922, `RNS_PRIME_BITS'd1590975914, `RNS_PRIME_BITS'd1400398196, `RNS_PRIME_BITS'd1787450196, `RNS_PRIME_BITS'd1560206244, `RNS_PRIME_BITS'd1107439066, `RNS_PRIME_BITS'd939528947, `RNS_PRIME_BITS'd1968363549},
    '{`RNS_PRIME_BITS'd110, `RNS_PRIME_BITS'd1259738977, `RNS_PRIME_BITS'd661307223, `RNS_PRIME_BITS'd1471575600, `RNS_PRIME_BITS'd1224673918, `RNS_PRIME_BITS'd782037768, `RNS_PRIME_BITS'd1168354671, `RNS_PRIME_BITS'd1705579202, `RNS_PRIME_BITS'd2041561652, `RNS_PRIME_BITS'd412736448, `RNS_PRIME_BITS'd1797787298},
    '{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd529873326, `RNS_PRIME_BITS'd1643627778, `RNS_PRIME_BITS'd176640802, `RNS_PRIME_BITS'd800805372, `RNS_PRIME_BITS'd2079567620, `RNS_PRIME_BITS'd1634430713, `RNS_PRIME_BITS'd381351274, `RNS_PRIME_BITS'd84392424, `RNS_PRIME_BITS'd1907477980, `RNS_PRIME_BITS'd173024403},
    '{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd1798433420, `RNS_PRIME_BITS'd426691550, `RNS_PRIME_BITS'd2046591696, `RNS_PRIME_BITS'd1896915698, `RNS_PRIME_BITS'd1668408377, `RNS_PRIME_BITS'd1455614987, `RNS_PRIME_BITS'd122326003, `RNS_PRIME_BITS'd298471715, `RNS_PRIME_BITS'd988993182, `RNS_PRIME_BITS'd973820226},
    '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1746944147, `RNS_PRIME_BITS'd689413926, `RNS_PRIME_BITS'd568471330, `RNS_PRIME_BITS'd236800200, `RNS_PRIME_BITS'd122139163, `RNS_PRIME_BITS'd1844962837, `RNS_PRIME_BITS'd2046340205, `RNS_PRIME_BITS'd1752607833, `RNS_PRIME_BITS'd38992541, `RNS_PRIME_BITS'd666891990},
    '{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd780035198, `RNS_PRIME_BITS'd696210963, `RNS_PRIME_BITS'd2088411844, `RNS_PRIME_BITS'd1803926386, `RNS_PRIME_BITS'd1141553323, `RNS_PRIME_BITS'd857805866, `RNS_PRIME_BITS'd460171280, `RNS_PRIME_BITS'd1285011956, `RNS_PRIME_BITS'd398309668, `RNS_PRIME_BITS'd1149897307},
    '{`RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd187755373, `RNS_PRIME_BITS'd290063258, `RNS_PRIME_BITS'd144189587, `RNS_PRIME_BITS'd264727076, `RNS_PRIME_BITS'd1186399849, `RNS_PRIME_BITS'd1391700885, `RNS_PRIME_BITS'd475214179, `RNS_PRIME_BITS'd103801546, `RNS_PRIME_BITS'd831416656, `RNS_PRIME_BITS'd694183001},
    '{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd1504604024, `RNS_PRIME_BITS'd2051724077, `RNS_PRIME_BITS'd460984520, `RNS_PRIME_BITS'd505776640, `RNS_PRIME_BITS'd1257572391, `RNS_PRIME_BITS'd619517657, `RNS_PRIME_BITS'd1520366584, `RNS_PRIME_BITS'd588667643, `RNS_PRIME_BITS'd613176604, `RNS_PRIME_BITS'd1678891938},
    '{`RNS_PRIME_BITS'd204, `RNS_PRIME_BITS'd87626930, `RNS_PRIME_BITS'd1428342435, `RNS_PRIME_BITS'd334829787, `RNS_PRIME_BITS'd575426957, `RNS_PRIME_BITS'd1135762866, `RNS_PRIME_BITS'd2028759844, `RNS_PRIME_BITS'd1925903783, `RNS_PRIME_BITS'd1137575117, `RNS_PRIME_BITS'd2035276103, `RNS_PRIME_BITS'd752620199},
    '{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd1472894111, `RNS_PRIME_BITS'd666024267, `RNS_PRIME_BITS'd161246845, `RNS_PRIME_BITS'd770546543, `RNS_PRIME_BITS'd264543334, `RNS_PRIME_BITS'd1156921900, `RNS_PRIME_BITS'd347183033, `RNS_PRIME_BITS'd1952749081, `RNS_PRIME_BITS'd135120200, `RNS_PRIME_BITS'd816699827}
};

`endif