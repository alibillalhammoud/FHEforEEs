`ifndef TYPES_SVH
`define TYPES_SVH

// ---------------------------
// Basic data types
// ---------------------------



// NTT
`define BASE      32'd2
// Width of each RNS residue (one small prime)
`define RNS_PRIME_BITS 32
// RNS residues
typedef logic [`RNS_PRIME_BITS-1:0] rns_residue_t; 
typedef logic [(2*`RNS_PRIME_BITS)-1:0] wide_rns_residue_t;
// Vector / slot params
`define N_SLOTS   64
// moduli and RNS bases
`define t_MODULUS 257

`define q_BASIS_LEN 11
//`define q_MODULUS = 536092687689737712660299305370020840707037344303743567681198293980556215074372863278673727266177
parameter rns_residue_t q_BASIS [`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353};
//`define B_MODULUS = 2086045702160390514072457421164142647843268814746900546792219301529141418454085790414389880321
`define B_BASIS_LEN 10
parameter rns_residue_t B_BASIS [`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337};
//`define Ba_MODULUS = 2147503489
`define Ba_BASIS_LEN 1
parameter rns_residue_t Ba_BASIS [`Ba_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147503489};
`define qBBa_BASIS_LEN 22
//`define qBBa_MODULUS = 2401582888476023779443294070753805757615044045174800139284098902756577490274881128570727198734820745298450301532339857214864378319647024214690248526201090429246246041638715397173165827069546764128513
parameter rns_residue_t qBBa_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353, `RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147503489};

parameter rns_residue_t w_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1684230034, `RNS_PRIME_BITS'd413528229, `RNS_PRIME_BITS'd835068854, `RNS_PRIME_BITS'd698897645, `RNS_PRIME_BITS'd266488565, `RNS_PRIME_BITS'd1915797300, `RNS_PRIME_BITS'd634442553, `RNS_PRIME_BITS'd207695132, `RNS_PRIME_BITS'd21725588, `RNS_PRIME_BITS'd209219715, `RNS_PRIME_BITS'd1654849230, `RNS_PRIME_BITS'd318222520, `RNS_PRIME_BITS'd458644985, `RNS_PRIME_BITS'd1659477478, `RNS_PRIME_BITS'd221897449, `RNS_PRIME_BITS'd1817702166, `RNS_PRIME_BITS'd1453892451, `RNS_PRIME_BITS'd1033346514, `RNS_PRIME_BITS'd1445995283, `RNS_PRIME_BITS'd330138710, `RNS_PRIME_BITS'd545722081};
parameter rns_residue_t w_INV_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd165, `RNS_PRIME_BITS'd465883484, `RNS_PRIME_BITS'd1309966555, `RNS_PRIME_BITS'd1089826325, `RNS_PRIME_BITS'd123767386, `RNS_PRIME_BITS'd1570352642, `RNS_PRIME_BITS'd374598187, `RNS_PRIME_BITS'd199676388, `RNS_PRIME_BITS'd1965833606, `RNS_PRIME_BITS'd1344902099, `RNS_PRIME_BITS'd1350503019, `RNS_PRIME_BITS'd1320961193, `RNS_PRIME_BITS'd1595145660, `RNS_PRIME_BITS'd673021473, `RNS_PRIME_BITS'd1565830187, `RNS_PRIME_BITS'd46526017, `RNS_PRIME_BITS'd1553448153, `RNS_PRIME_BITS'd1394618113, `RNS_PRIME_BITS'd1852124673, `RNS_PRIME_BITS'd1285194286, `RNS_PRIME_BITS'd438577756, `RNS_PRIME_BITS'd433881419};

`define BBa_BASIS_LEN 11
parameter rns_residue_t BBa_BASIS [`BBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147503489};

// RNS integers
typedef rns_residue_t rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef rns_residue_t rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef rns_residue_t rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
typedef rns_residue_t rns_coef_qBBa_BASIS_t [`q_BASIS_LEN + `B_BASIS_LEN + `Ba_BASIS_LEN];
typedef rns_residue_t rns_coef_BBa_BASIS_t [`B_BASIS_LEN + `Ba_BASIS_LEN];
// Polynomials
typedef rns_int_q_BASIS_t q_BASIS_poly [`N_SLOTS]; 
typedef rns_int_B_BASIS_t B_BASIS_poly [`N_SLOTS]; 
typedef rns_int_Ba_BASIS_t Ba_BASIS_poly [`N_SLOTS];
typedef rns_coef_BBa_BASIS_t BBa_BASIS_poly [`N_SLOTS];
typedef rns_coef_qBBa_BASIS_t qBBa_BASIS_poly [`N_SLOTS];
// wide RNS integers (each residue is double the length for mult)
typedef wide_rns_residue_t wide_rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
// wide Polynomials
typedef wide_rns_int_q_BASIS_t wide_q_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_B_BASIS_t wide_B_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_Ba_BASIS_t wide_Ba_BASIS_poly [`N_SLOTS];

// ---------------------------
// precalculated values
// ---------------------------
// NTT precalculated factors

// parameter q_BASIS_poly twist_factor_q = '{default: 1'b1};
// parameter B_BASIS_poly twist_factor_b = '{default: 1'b1};
// parameter Ba_BASIS_poly twist_factor_ba = '{default: 1'b1};

// parameter q_BASIS_poly untwist_factor_q = '{default: 1'b1};
// parameter b_BASIS_poly untwist_factor_b = '{default: 1'b1};
// parameter q_BASIS_poly untwist_factor_ba = '{default: 1'b1};


parameter q_BASIS_poly twist_factor_q   = '{
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1},
    '{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1454056114, `RNS_PRIME_BITS'd2023476074, `RNS_PRIME_BITS'd1829761212, `RNS_PRIME_BITS'd1180811958, `RNS_PRIME_BITS'd863581131, `RNS_PRIME_BITS'd2006888302, `RNS_PRIME_BITS'd827630191, `RNS_PRIME_BITS'd1925970851, `RNS_PRIME_BITS'd679082962, `RNS_PRIME_BITS'd985627742},
    '{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1684230034, `RNS_PRIME_BITS'd413528229, `RNS_PRIME_BITS'd835068854, `RNS_PRIME_BITS'd698897645, `RNS_PRIME_BITS'd266488565, `RNS_PRIME_BITS'd1915797300, `RNS_PRIME_BITS'd634442553, `RNS_PRIME_BITS'd207695132, `RNS_PRIME_BITS'd21725588, `RNS_PRIME_BITS'd209219715},
    '{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd1874017521, `RNS_PRIME_BITS'd1276327416, `RNS_PRIME_BITS'd765723923, `RNS_PRIME_BITS'd396752410, `RNS_PRIME_BITS'd197474481, `RNS_PRIME_BITS'd49249814, `RNS_PRIME_BITS'd14124402, `RNS_PRIME_BITS'd148848534, `RNS_PRIME_BITS'd1645223958, `RNS_PRIME_BITS'd1797297359},
    '{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd120548658, `RNS_PRIME_BITS'd67511054, `RNS_PRIME_BITS'd346940440, `RNS_PRIME_BITS'd1590960824, `RNS_PRIME_BITS'd2131754249, `RNS_PRIME_BITS'd1610378484, `RNS_PRIME_BITS'd1687474151, `RNS_PRIME_BITS'd1761745303, `RNS_PRIME_BITS'd1935386753, `RNS_PRIME_BITS'd607947504},
    '{`RNS_PRIME_BITS'd196, `RNS_PRIME_BITS'd340182173, `RNS_PRIME_BITS'd951629099, `RNS_PRIME_BITS'd538002895, `RNS_PRIME_BITS'd676858767, `RNS_PRIME_BITS'd1844273609, `RNS_PRIME_BITS'd808269908, `RNS_PRIME_BITS'd14861374, `RNS_PRIME_BITS'd1020094163, `RNS_PRIME_BITS'd147309818, `RNS_PRIME_BITS'd582137866},
    '{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd656530581, `RNS_PRIME_BITS'd861227005, `RNS_PRIME_BITS'd1064440654, `RNS_PRIME_BITS'd1242864821, `RNS_PRIME_BITS'd2052452190, `RNS_PRIME_BITS'd1579153117, `RNS_PRIME_BITS'd1248849378, `RNS_PRIME_BITS'd1296504500, `RNS_PRIME_BITS'd1358855180, `RNS_PRIME_BITS'd1553772574},
    '{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd1079385897, `RNS_PRIME_BITS'd576378926, `RNS_PRIME_BITS'd1614098500, `RNS_PRIME_BITS'd1981568237, `RNS_PRIME_BITS'd1532049341, `RNS_PRIME_BITS'd785126063, `RNS_PRIME_BITS'd2105098028, `RNS_PRIME_BITS'd1590156063, `RNS_PRIME_BITS'd1309811091, `RNS_PRIME_BITS'd1001224375},
    '{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd1323801281, `RNS_PRIME_BITS'd1485798473, `RNS_PRIME_BITS'd469931230, `RNS_PRIME_BITS'd2047801397, `RNS_PRIME_BITS'd1811004807, `RNS_PRIME_BITS'd1519044505, `RNS_PRIME_BITS'd1655854283, `RNS_PRIME_BITS'd1828920336, `RNS_PRIME_BITS'd1178694670, `RNS_PRIME_BITS'd408115440},
    '{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd1753733667, `RNS_PRIME_BITS'd857515399, `RNS_PRIME_BITS'd1345302327, `RNS_PRIME_BITS'd1141109968, `RNS_PRIME_BITS'd1970163605, `RNS_PRIME_BITS'd1343154438, `RNS_PRIME_BITS'd1376784415, `RNS_PRIME_BITS'd1528595831, `RNS_PRIME_BITS'd1626480704, `RNS_PRIME_BITS'd1688164042},
    '{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd109329595, `RNS_PRIME_BITS'd1603393679, `RNS_PRIME_BITS'd1699086710, `RNS_PRIME_BITS'd640452388, `RNS_PRIME_BITS'd1802277828, `RNS_PRIME_BITS'd106304448, `RNS_PRIME_BITS'd1875735111, `RNS_PRIME_BITS'd1612223517, `RNS_PRIME_BITS'd789699425, `RNS_PRIME_BITS'd1138957206},
    '{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1102767568, `RNS_PRIME_BITS'd1804390941, `RNS_PRIME_BITS'd190235933, `RNS_PRIME_BITS'd1735615176, `RNS_PRIME_BITS'd200129577, `RNS_PRIME_BITS'd1361590782, `RNS_PRIME_BITS'd1629799445, `RNS_PRIME_BITS'd1146443053, `RNS_PRIME_BITS'd1362151287, `RNS_PRIME_BITS'd29488642},
    '{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd2066618854, `RNS_PRIME_BITS'd1867409965, `RNS_PRIME_BITS'd973917268, `RNS_PRIME_BITS'd104371406, `RNS_PRIME_BITS'd1902288884, `RNS_PRIME_BITS'd408243051, `RNS_PRIME_BITS'd50859102, `RNS_PRIME_BITS'd822124619, `RNS_PRIME_BITS'd1335637725, `RNS_PRIME_BITS'd695959640},
    '{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd1323556320, `RNS_PRIME_BITS'd2064658918, `RNS_PRIME_BITS'd1573977587, `RNS_PRIME_BITS'd793743842, `RNS_PRIME_BITS'd600242329, `RNS_PRIME_BITS'd1624358720, `RNS_PRIME_BITS'd353092123, `RNS_PRIME_BITS'd373441180, `RNS_PRIME_BITS'd799792040, `RNS_PRIME_BITS'd1479303328},
    '{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd668212887, `RNS_PRIME_BITS'd1957088536, `RNS_PRIME_BITS'd765942372, `RNS_PRIME_BITS'd1404190271, `RNS_PRIME_BITS'd400413469, `RNS_PRIME_BITS'd1076916254, `RNS_PRIME_BITS'd1463329648, `RNS_PRIME_BITS'd1599886708, `RNS_PRIME_BITS'd1787703015, `RNS_PRIME_BITS'd519154132},
    '{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1871724384, `RNS_PRIME_BITS'd1016906757, `RNS_PRIME_BITS'd631590787, `RNS_PRIME_BITS'd404036694, `RNS_PRIME_BITS'd735419640, `RNS_PRIME_BITS'd1411883997, `RNS_PRIME_BITS'd1971964208, `RNS_PRIME_BITS'd1819024442, `RNS_PRIME_BITS'd1889383441, `RNS_PRIME_BITS'd963399678},
    '{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd1061363846, `RNS_PRIME_BITS'd2093569547, `RNS_PRIME_BITS'd239311507, `RNS_PRIME_BITS'd2100155542, `RNS_PRIME_BITS'd10234283, `RNS_PRIME_BITS'd1499897549, `RNS_PRIME_BITS'd1351991644, `RNS_PRIME_BITS'd1343916693, `RNS_PRIME_BITS'd376392512, `RNS_PRIME_BITS'd405602459},
    '{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd248740266, `RNS_PRIME_BITS'd1953159839, `RNS_PRIME_BITS'd793606413, `RNS_PRIME_BITS'd1947317042, `RNS_PRIME_BITS'd1236975143, `RNS_PRIME_BITS'd995275098, `RNS_PRIME_BITS'd1423704554, `RNS_PRIME_BITS'd1580226385, `RNS_PRIME_BITS'd1203126727, `RNS_PRIME_BITS'd1892086515},
    '{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd918758775, `RNS_PRIME_BITS'd74609970, `RNS_PRIME_BITS'd1368161792, `RNS_PRIME_BITS'd1002584402, `RNS_PRIME_BITS'd354809650, `RNS_PRIME_BITS'd573382855, `RNS_PRIME_BITS'd462906762, `RNS_PRIME_BITS'd1465397025, `RNS_PRIME_BITS'd649865995, `RNS_PRIME_BITS'd80644722},
    '{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd1340620076, `RNS_PRIME_BITS'd435782459, `RNS_PRIME_BITS'd1256631702, `RNS_PRIME_BITS'd1972104903, `RNS_PRIME_BITS'd1260290827, `RNS_PRIME_BITS'd796043708, `RNS_PRIME_BITS'd1662891139, `RNS_PRIME_BITS'd576340174, `RNS_PRIME_BITS'd1898940369, `RNS_PRIME_BITS'd1766908121},
    '{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd1215568715, `RNS_PRIME_BITS'd764376413, `RNS_PRIME_BITS'd1968585711, `RNS_PRIME_BITS'd1117302355, `RNS_PRIME_BITS'd240751673, `RNS_PRIME_BITS'd1898906447, `RNS_PRIME_BITS'd1537383243, `RNS_PRIME_BITS'd508007782, `RNS_PRIME_BITS'd1306763942, `RNS_PRIME_BITS'd589212064},
    '{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd16030913, `RNS_PRIME_BITS'd1073050120, `RNS_PRIME_BITS'd56850842, `RNS_PRIME_BITS'd1082672190, `RNS_PRIME_BITS'd2076469305, `RNS_PRIME_BITS'd2046261189, `RNS_PRIME_BITS'd190823532, `RNS_PRIME_BITS'd1949278380, `RNS_PRIME_BITS'd896631706, `RNS_PRIME_BITS'd1938421324},
    '{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd1583075798, `RNS_PRIME_BITS'd599521406, `RNS_PRIME_BITS'd2122922145, `RNS_PRIME_BITS'd665909595, `RNS_PRIME_BITS'd231305546, `RNS_PRIME_BITS'd1898694097, `RNS_PRIME_BITS'd754518586, `RNS_PRIME_BITS'd1026065501, `RNS_PRIME_BITS'd1233985319, `RNS_PRIME_BITS'd223488580},
    '{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd702020947, `RNS_PRIME_BITS'd1695639893, `RNS_PRIME_BITS'd1904384299, `RNS_PRIME_BITS'd325883975, `RNS_PRIME_BITS'd122535444, `RNS_PRIME_BITS'd1866665936, `RNS_PRIME_BITS'd1472669913, `RNS_PRIME_BITS'd1982388385, `RNS_PRIME_BITS'd1297846148, `RNS_PRIME_BITS'd1007863781},
    '{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd426187835, `RNS_PRIME_BITS'd1884145470, `RNS_PRIME_BITS'd514016804, `RNS_PRIME_BITS'd1855667154, `RNS_PRIME_BITS'd1634152440, `RNS_PRIME_BITS'd321460536, `RNS_PRIME_BITS'd1403908978, `RNS_PRIME_BITS'd601571399, `RNS_PRIME_BITS'd1971934677, `RNS_PRIME_BITS'd572067441},
    '{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1577612670, `RNS_PRIME_BITS'd1387757027, `RNS_PRIME_BITS'd1634409210, `RNS_PRIME_BITS'd536371151, `RNS_PRIME_BITS'd449910378, `RNS_PRIME_BITS'd1935227906, `RNS_PRIME_BITS'd838777520, `RNS_PRIME_BITS'd1814968618, `RNS_PRIME_BITS'd1424335466, `RNS_PRIME_BITS'd1628177047},
    '{`RNS_PRIME_BITS'd162, `RNS_PRIME_BITS'd994527522, `RNS_PRIME_BITS'd837323404, `RNS_PRIME_BITS'd552952089, `RNS_PRIME_BITS'd431097772, `RNS_PRIME_BITS'd1239381293, `RNS_PRIME_BITS'd292174375, `RNS_PRIME_BITS'd356624563, `RNS_PRIME_BITS'd1139796275, `RNS_PRIME_BITS'd216329546, `RNS_PRIME_BITS'd70232036},
    '{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd994513885, `RNS_PRIME_BITS'd1449362922, `RNS_PRIME_BITS'd257231880, `RNS_PRIME_BITS'd1527060402, `RNS_PRIME_BITS'd2113046598, `RNS_PRIME_BITS'd1651256030, `RNS_PRIME_BITS'd1854365554, `RNS_PRIME_BITS'd1376844757, `RNS_PRIME_BITS'd1938315192, `RNS_PRIME_BITS'd888471290},
    '{`RNS_PRIME_BITS'd15, `RNS_PRIME_BITS'd1896484085, `RNS_PRIME_BITS'd1456040658, `RNS_PRIME_BITS'd998069335, `RNS_PRIME_BITS'd1113343725, `RNS_PRIME_BITS'd1065183214, `RNS_PRIME_BITS'd1674111577, `RNS_PRIME_BITS'd1405622643, `RNS_PRIME_BITS'd591326689, `RNS_PRIME_BITS'd1163148101, `RNS_PRIME_BITS'd41854895},
    '{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd1390505442, `RNS_PRIME_BITS'd1703996997, `RNS_PRIME_BITS'd132272763, `RNS_PRIME_BITS'd1952670695, `RNS_PRIME_BITS'd523000083, `RNS_PRIME_BITS'd362735615, `RNS_PRIME_BITS'd182689866, `RNS_PRIME_BITS'd284129690, `RNS_PRIME_BITS'd1843731486, `RNS_PRIME_BITS'd369428266},
    '{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd470517865, `RNS_PRIME_BITS'd1343049929, `RNS_PRIME_BITS'd242912769, `RNS_PRIME_BITS'd1494908283, `RNS_PRIME_BITS'd831666628, `RNS_PRIME_BITS'd303641034, `RNS_PRIME_BITS'd2088866633, `RNS_PRIME_BITS'd1468519535, `RNS_PRIME_BITS'd2000376334, `RNS_PRIME_BITS'd980564471},
    '{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd1521041901, `RNS_PRIME_BITS'd788800085, `RNS_PRIME_BITS'd185065907, `RNS_PRIME_BITS'd1889283537, `RNS_PRIME_BITS'd138524561, `RNS_PRIME_BITS'd136679130, `RNS_PRIME_BITS'd1993147357, `RNS_PRIME_BITS'd827950938, `RNS_PRIME_BITS'd153601635, `RNS_PRIME_BITS'd1490691155},
    '{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd1021707020, `RNS_PRIME_BITS'd434575099, `RNS_PRIME_BITS'd1712127733, `RNS_PRIME_BITS'd524962442, `RNS_PRIME_BITS'd1172437812, `RNS_PRIME_BITS'd947974746, `RNS_PRIME_BITS'd335862598, `RNS_PRIME_BITS'd1331495236, `RNS_PRIME_BITS'd1410137926, `RNS_PRIME_BITS'd37028611},
    '{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd774040236, `RNS_PRIME_BITS'd572591813, `RNS_PRIME_BITS'd1210603202, `RNS_PRIME_BITS'd1401061297, `RNS_PRIME_BITS'd590795774, `RNS_PRIME_BITS'd1971088069, `RNS_PRIME_BITS'd520746293, `RNS_PRIME_BITS'd1575358450, `RNS_PRIME_BITS'd476307234, `RNS_PRIME_BITS'd2016849603},
    '{`RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd42370405, `RNS_PRIME_BITS'd813012214, `RNS_PRIME_BITS'd1479849359, `RNS_PRIME_BITS'd1349253646, `RNS_PRIME_BITS'd348980417, `RNS_PRIME_BITS'd331719264, `RNS_PRIME_BITS'd795266135, `RNS_PRIME_BITS'd368435717, `RNS_PRIME_BITS'd489843704, `RNS_PRIME_BITS'd269448364},
    '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1260414647, `RNS_PRIME_BITS'd1319821704, `RNS_PRIME_BITS'd618256455, `RNS_PRIME_BITS'd818503666, `RNS_PRIME_BITS'd1897963711, `RNS_PRIME_BITS'd1067104690, `RNS_PRIME_BITS'd276444971, `RNS_PRIME_BITS'd1380291710, `RNS_PRIME_BITS'd1154289721, `RNS_PRIME_BITS'd1080531861},
    '{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd2121222217, `RNS_PRIME_BITS'd1458297369, `RNS_PRIME_BITS'd336159836, `RNS_PRIME_BITS'd723680490, `RNS_PRIME_BITS'd1718005309, `RNS_PRIME_BITS'd1014920853, `RNS_PRIME_BITS'd1008493454, `RNS_PRIME_BITS'd353025982, `RNS_PRIME_BITS'd741963136, `RNS_PRIME_BITS'd117506787},
    '{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd1547276440, `RNS_PRIME_BITS'd688415855, `RNS_PRIME_BITS'd618238460, `RNS_PRIME_BITS'd322476241, `RNS_PRIME_BITS'd1133296249, `RNS_PRIME_BITS'd447649351, `RNS_PRIME_BITS'd1962983607, `RNS_PRIME_BITS'd228998489, `RNS_PRIME_BITS'd205108911, `RNS_PRIME_BITS'd1446317206},
    '{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd1934841955, `RNS_PRIME_BITS'd34272266, `RNS_PRIME_BITS'd1169566253, `RNS_PRIME_BITS'd1874038872, `RNS_PRIME_BITS'd796514801, `RNS_PRIME_BITS'd305771017, `RNS_PRIME_BITS'd737870517, `RNS_PRIME_BITS'd1188901935, `RNS_PRIME_BITS'd1051329728, `RNS_PRIME_BITS'd1362925816},
    '{`RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd883135528, `RNS_PRIME_BITS'd514568416, `RNS_PRIME_BITS'd1653743872, `RNS_PRIME_BITS'd834025286, `RNS_PRIME_BITS'd958676669, `RNS_PRIME_BITS'd959695467, `RNS_PRIME_BITS'd140078324, `RNS_PRIME_BITS'd1389915387, `RNS_PRIME_BITS'd881212437, `RNS_PRIME_BITS'd702116429},
    '{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1146745373, `RNS_PRIME_BITS'd108956348, `RNS_PRIME_BITS'd230876332, `RNS_PRIME_BITS'd281055234, `RNS_PRIME_BITS'd64563004, `RNS_PRIME_BITS'd731192465, `RNS_PRIME_BITS'd608663139, `RNS_PRIME_BITS'd464898846, `RNS_PRIME_BITS'd1454002446, `RNS_PRIME_BITS'd1232945780},
    '{`RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd501271165, `RNS_PRIME_BITS'd1695216211, `RNS_PRIME_BITS'd1199214675, `RNS_PRIME_BITS'd1074140584, `RNS_PRIME_BITS'd1975647812, `RNS_PRIME_BITS'd596300382, `RNS_PRIME_BITS'd481530671, `RNS_PRIME_BITS'd1250107969, `RNS_PRIME_BITS'd59717368, `RNS_PRIME_BITS'd410918689},
    '{`RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd788019979, `RNS_PRIME_BITS'd1530978778, `RNS_PRIME_BITS'd1878325668, `RNS_PRIME_BITS'd49981851, `RNS_PRIME_BITS'd579138741, `RNS_PRIME_BITS'd1769119785, `RNS_PRIME_BITS'd1794412482, `RNS_PRIME_BITS'd622888137, `RNS_PRIME_BITS'd1546369699, `RNS_PRIME_BITS'd156420353},
    '{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd1009909057, `RNS_PRIME_BITS'd1563397195, `RNS_PRIME_BITS'd7727696, `RNS_PRIME_BITS'd878592647, `RNS_PRIME_BITS'd36175035, `RNS_PRIME_BITS'd1902426573, `RNS_PRIME_BITS'd944136518, `RNS_PRIME_BITS'd87729872, `RNS_PRIME_BITS'd1009475440, `RNS_PRIME_BITS'd901760470},
    '{`RNS_PRIME_BITS'd189, `RNS_PRIME_BITS'd1963269275, `RNS_PRIME_BITS'd1871639102, `RNS_PRIME_BITS'd909482893, `RNS_PRIME_BITS'd1280361918, `RNS_PRIME_BITS'd182951808, `RNS_PRIME_BITS'd654833583, `RNS_PRIME_BITS'd1479984746, `RNS_PRIME_BITS'd1083576085, `RNS_PRIME_BITS'd539509008, `RNS_PRIME_BITS'd1589572379},
    '{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd1270209618, `RNS_PRIME_BITS'd572522453, `RNS_PRIME_BITS'd390894248, `RNS_PRIME_BITS'd1657938546, `RNS_PRIME_BITS'd1491813251, `RNS_PRIME_BITS'd873629554, `RNS_PRIME_BITS'd1020523066, `RNS_PRIME_BITS'd1840014191, `RNS_PRIME_BITS'd341138130, `RNS_PRIME_BITS'd472182866},
    '{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd763626807, `RNS_PRIME_BITS'd1339861729, `RNS_PRIME_BITS'd791713145, `RNS_PRIME_BITS'd658448763, `RNS_PRIME_BITS'd1193767449, `RNS_PRIME_BITS'd711101770, `RNS_PRIME_BITS'd1308174171, `RNS_PRIME_BITS'd1453536448, `RNS_PRIME_BITS'd1720619438, `RNS_PRIME_BITS'd1578477615},
    '{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd480335015, `RNS_PRIME_BITS'd800312580, `RNS_PRIME_BITS'd1215966900, `RNS_PRIME_BITS'd1234006662, `RNS_PRIME_BITS'd1756567829, `RNS_PRIME_BITS'd679149815, `RNS_PRIME_BITS'd129364822, `RNS_PRIME_BITS'd1893528272, `RNS_PRIME_BITS'd535596838, `RNS_PRIME_BITS'd1370829515},
    '{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd910119688, `RNS_PRIME_BITS'd1128292512, `RNS_PRIME_BITS'd587075636, `RNS_PRIME_BITS'd1800184525, `RNS_PRIME_BITS'd1221476635, `RNS_PRIME_BITS'd558407411, `RNS_PRIME_BITS'd1843702908, `RNS_PRIME_BITS'd824257829, `RNS_PRIME_BITS'd1631833303, `RNS_PRIME_BITS'd2028194232},
    '{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1159872543, `RNS_PRIME_BITS'd1784665556, `RNS_PRIME_BITS'd1199234809, `RNS_PRIME_BITS'd1599760116, `RNS_PRIME_BITS'd1663696998, `RNS_PRIME_BITS'd449470596, `RNS_PRIME_BITS'd1806730708, `RNS_PRIME_BITS'd923463583, `RNS_PRIME_BITS'd933766656, `RNS_PRIME_BITS'd971006858},
    '{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd1182896170, `RNS_PRIME_BITS'd113138122, `RNS_PRIME_BITS'd39126152, `RNS_PRIME_BITS'd1944520926, `RNS_PRIME_BITS'd1660937547, `RNS_PRIME_BITS'd276205002, `RNS_PRIME_BITS'd688071846, `RNS_PRIME_BITS'd1538410082, `RNS_PRIME_BITS'd926729148, `RNS_PRIME_BITS'd908554640},
    '{`RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd350490837, `RNS_PRIME_BITS'd228923992, `RNS_PRIME_BITS'd624524991, `RNS_PRIME_BITS'd1201959893, `RNS_PRIME_BITS'd19608843, `RNS_PRIME_BITS'd1788733215, `RNS_PRIME_BITS'd2031608751, `RNS_PRIME_BITS'd1174453731, `RNS_PRIME_BITS'd1837590264, `RNS_PRIME_BITS'd768568972},
    '{`RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd2086471810, `RNS_PRIME_BITS'd31790164, `RNS_PRIME_BITS'd1200643284, `RNS_PRIME_BITS'd1601517741, `RNS_PRIME_BITS'd1804134098, `RNS_PRIME_BITS'd429865127, `RNS_PRIME_BITS'd1141675715, `RNS_PRIME_BITS'd911258653, `RNS_PRIME_BITS'd621781956, `RNS_PRIME_BITS'd202469597},
    '{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd1074706051, `RNS_PRIME_BITS'd183046999, `RNS_PRIME_BITS'd2068724100, `RNS_PRIME_BITS'd366288311, `RNS_PRIME_BITS'd1143024219, `RNS_PRIME_BITS'd1275811230, `RNS_PRIME_BITS'd2018762224, `RNS_PRIME_BITS'd712118336, `RNS_PRIME_BITS'd2122931229, `RNS_PRIME_BITS'd1343706043},
    '{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd248908061, `RNS_PRIME_BITS'd984227194, `RNS_PRIME_BITS'd1028019199, `RNS_PRIME_BITS'd1067917992, `RNS_PRIME_BITS'd887687435, `RNS_PRIME_BITS'd1370277766, `RNS_PRIME_BITS'd999896244, `RNS_PRIME_BITS'd1078820638, `RNS_PRIME_BITS'd2098610929, `RNS_PRIME_BITS'd387366877},
    '{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd42567327, `RNS_PRIME_BITS'd1940067462, `RNS_PRIME_BITS'd764503116, `RNS_PRIME_BITS'd1471009666, `RNS_PRIME_BITS'd1287398144, `RNS_PRIME_BITS'd1168169987, `RNS_PRIME_BITS'd703901652, `RNS_PRIME_BITS'd1901471095, `RNS_PRIME_BITS'd863275331, `RNS_PRIME_BITS'd1612097702},
    '{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd1605683, `RNS_PRIME_BITS'd397906100, `RNS_PRIME_BITS'd956844079, `RNS_PRIME_BITS'd1724844730, `RNS_PRIME_BITS'd120671020, `RNS_PRIME_BITS'd538488167, `RNS_PRIME_BITS'd1469183668, `RNS_PRIME_BITS'd768800080, `RNS_PRIME_BITS'd1075515373, `RNS_PRIME_BITS'd316054804},
    '{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd231006354, `RNS_PRIME_BITS'd377036607, `RNS_PRIME_BITS'd976022455, `RNS_PRIME_BITS'd1186389507, `RNS_PRIME_BITS'd660093495, `RNS_PRIME_BITS'd126138005, `RNS_PRIME_BITS'd1633319106, `RNS_PRIME_BITS'd1427536931, `RNS_PRIME_BITS'd375638505, `RNS_PRIME_BITS'd400914411},
    '{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd328404460, `RNS_PRIME_BITS'd1578585534, `RNS_PRIME_BITS'd128768493, `RNS_PRIME_BITS'd1232517567, `RNS_PRIME_BITS'd1773444005, `RNS_PRIME_BITS'd1843645976, `RNS_PRIME_BITS'd541653944, `RNS_PRIME_BITS'd1721350193, `RNS_PRIME_BITS'd665726026, `RNS_PRIME_BITS'd828730173},
    '{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd184517896, `RNS_PRIME_BITS'd1760756591, `RNS_PRIME_BITS'd601425161, `RNS_PRIME_BITS'd2054892602, `RNS_PRIME_BITS'd960444154, `RNS_PRIME_BITS'd342817420, `RNS_PRIME_BITS'd1165857483, `RNS_PRIME_BITS'd421031535, `RNS_PRIME_BITS'd467316107, `RNS_PRIME_BITS'd786533504},
    '{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd1628067296, `RNS_PRIME_BITS'd445410876, `RNS_PRIME_BITS'd297804970, `RNS_PRIME_BITS'd1556827466, `RNS_PRIME_BITS'd1827198507, `RNS_PRIME_BITS'd667896261, `RNS_PRIME_BITS'd187415820, `RNS_PRIME_BITS'd1756461716, `RNS_PRIME_BITS'd547754318, `RNS_PRIME_BITS'd574179569},
    '{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd1495990324, `RNS_PRIME_BITS'd384884134, `RNS_PRIME_BITS'd86626384, `RNS_PRIME_BITS'd971038417, `RNS_PRIME_BITS'd1783905120, `RNS_PRIME_BITS'd1326718868, `RNS_PRIME_BITS'd1347391675, `RNS_PRIME_BITS'd1423546356, `RNS_PRIME_BITS'd1580566206, `RNS_PRIME_BITS'd935110882},
    '{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd1681600293, `RNS_PRIME_BITS'd837517606, `RNS_PRIME_BITS'd1057658604, `RNS_PRIME_BITS'd2023717671, `RNS_PRIME_BITS'd577134207, `RNS_PRIME_BITS'd1772889814, `RNS_PRIME_BITS'd1947813149, `RNS_PRIME_BITS'd181657083, `RNS_PRIME_BITS'd802589102, `RNS_PRIME_BITS'd796989334},
    '{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1180703254, `RNS_PRIME_BITS'd718232802, `RNS_PRIME_BITS'd1158945815, `RNS_PRIME_BITS'd1674979427, `RNS_PRIME_BITS'd708871736, `RNS_PRIME_BITS'd1423092132, `RNS_PRIME_BITS'd1192713535, `RNS_PRIME_BITS'd1451070185, `RNS_PRIME_BITS'd148205767, `RNS_PRIME_BITS'd732343142}
};
parameter q_BASIS_poly untwist_factor_q = '{
    '{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd2113929343, `RNS_PRIME_BITS'd2113929721, `RNS_PRIME_BITS'd2113930477, `RNS_PRIME_BITS'd2113930603, `RNS_PRIME_BITS'd2113932367, `RNS_PRIME_BITS'd2113933501, `RNS_PRIME_BITS'd2113935013, `RNS_PRIME_BITS'd2113936147, `RNS_PRIME_BITS'd2113936651, `RNS_PRIME_BITS'd2113937785},
    '{`RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd719749060, `RNS_PRIME_BITS'd1129628573, `RNS_PRIME_BITS'd753643868, `RNS_PRIME_BITS'd1148234337, `RNS_PRIME_BITS'd1867974872, `RNS_PRIME_BITS'd1185726186, `RNS_PRIME_BITS'd2095298864, `RNS_PRIME_BITS'd1353063251, `RNS_PRIME_BITS'd232566135, `RNS_PRIME_BITS'd1263630723},
    '{`RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd1215239054, `RNS_PRIME_BITS'd1261982508, `RNS_PRIME_BITS'd1459869973, `RNS_PRIME_BITS'd1277003118, `RNS_PRIME_BITS'd2104914645, `RNS_PRIME_BITS'd710497597, `RNS_PRIME_BITS'd942646616, `RNS_PRIME_BITS'd1976879587, `RNS_PRIME_BITS'd1530968846, `RNS_PRIME_BITS'd725747538},
    '{`RNS_PRIME_BITS'd98, `RNS_PRIME_BITS'd1721455720, `RNS_PRIME_BITS'd1269054906, `RNS_PRIME_BITS'd535517695, `RNS_PRIME_BITS'd555253243, `RNS_PRIME_BITS'd1045869907, `RNS_PRIME_BITS'd650360018, `RNS_PRIME_BITS'd1958663922, `RNS_PRIME_BITS'd1722593273, `RNS_PRIME_BITS'd2055685754, `RNS_PRIME_BITS'd1126244205},
    '{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd1048303337, `RNS_PRIME_BITS'd2006306856, `RNS_PRIME_BITS'd1404633782, `RNS_PRIME_BITS'd311219111, `RNS_PRIME_BITS'd1414292750, `RNS_PRIME_BITS'd157336621, `RNS_PRIME_BITS'd399725916, `RNS_PRIME_BITS'd643646126, `RNS_PRIME_BITS'd461205039, `RNS_PRIME_BITS'd1635202277},
    '{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd265552380, `RNS_PRIME_BITS'd1549546859, `RNS_PRIME_BITS'd292592800, `RNS_PRIME_BITS'd1914050636, `RNS_PRIME_BITS'd1931153017, `RNS_PRIME_BITS'd397297478, `RNS_PRIME_BITS'd350883241, `RNS_PRIME_BITS'd1570484857, `RNS_PRIME_BITS'd361798236, `RNS_PRIME_BITS'd2135202767},
    '{`RNS_PRIME_BITS'd169, `RNS_PRIME_BITS'd1471263777, `RNS_PRIME_BITS'd2055709882, `RNS_PRIME_BITS'd1507938333, `RNS_PRIME_BITS'd2094672516, `RNS_PRIME_BITS'd1213805772, `RNS_PRIME_BITS'd776501032, `RNS_PRIME_BITS'd1870590002, `RNS_PRIME_BITS'd1617276462, `RNS_PRIME_BITS'd325143531, `RNS_PRIME_BITS'd2033879740},
    '{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd600370338, `RNS_PRIME_BITS'd2108038524, `RNS_PRIME_BITS'd1830244510, `RNS_PRIME_BITS'd82126026, `RNS_PRIME_BITS'd1835182550, `RNS_PRIME_BITS'd702673594, `RNS_PRIME_BITS'd41588437, `RNS_PRIME_BITS'd1152103706, `RNS_PRIME_BITS'd1369867199, `RNS_PRIME_BITS'd1436582137},
    '{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd1711251046, `RNS_PRIME_BITS'd1738613598, `RNS_PRIME_BITS'd1562108556, `RNS_PRIME_BITS'd1919207634, `RNS_PRIME_BITS'd1474511724, `RNS_PRIME_BITS'd1300211623, `RNS_PRIME_BITS'd1721879254, `RNS_PRIME_BITS'd524860171, `RNS_PRIME_BITS'd1493149823, `RNS_PRIME_BITS'd666153004},
    '{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd1039522340, `RNS_PRIME_BITS'd171013086, `RNS_PRIME_BITS'd390708063, `RNS_PRIME_BITS'd44124382, `RNS_PRIME_BITS'd2127371253, `RNS_PRIME_BITS'd82410844, `RNS_PRIME_BITS'd660092017, `RNS_PRIME_BITS'd1815789325, `RNS_PRIME_BITS'd87174973, `RNS_PRIME_BITS'd1249884558},
    '{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd969189398, `RNS_PRIME_BITS'd1930778971, `RNS_PRIME_BITS'd2097867677, `RNS_PRIME_BITS'd1325491942, `RNS_PRIME_BITS'd355229186, `RNS_PRIME_BITS'd179916410, `RNS_PRIME_BITS'd1729211870, `RNS_PRIME_BITS'd989779688, `RNS_PRIME_BITS'd1611382155, `RNS_PRIME_BITS'd967029865},
    '{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd83871020, `RNS_PRIME_BITS'd768892011, `RNS_PRIME_BITS'd101893994, `RNS_PRIME_BITS'd1839771716, `RNS_PRIME_BITS'd888111261, `RNS_PRIME_BITS'd986700450, `RNS_PRIME_BITS'd1579073993, `RNS_PRIME_BITS'd2136363840, `RNS_PRIME_BITS'd939911150, `RNS_PRIME_BITS'd1958724106},
    '{`RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd34507746, `RNS_PRIME_BITS'd670592079, `RNS_PRIME_BITS'd652328989, `RNS_PRIME_BITS'd1484926716, `RNS_PRIME_BITS'd575791081, `RNS_PRIME_BITS'd1301908858, `RNS_PRIME_BITS'd82824889, `RNS_PRIME_BITS'd958843302, `RNS_PRIME_BITS'd124502857, `RNS_PRIME_BITS'd969918885},
    '{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd699166695, `RNS_PRIME_BITS'd801729623, `RNS_PRIME_BITS'd2104172274, `RNS_PRIME_BITS'd685862911, `RNS_PRIME_BITS'd368792914, `RNS_PRIME_BITS'd1012240544, `RNS_PRIME_BITS'd1545318742, `RNS_PRIME_BITS'd1156058131, `RNS_PRIME_BITS'd1850342453, `RNS_PRIME_BITS'd390645926},
    '{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd1390803476, `RNS_PRIME_BITS'd333776617, `RNS_PRIME_BITS'd267824270, `RNS_PRIME_BITS'd976250481, `RNS_PRIME_BITS'd343147153, `RNS_PRIME_BITS'd331229297, `RNS_PRIME_BITS'd1264320790, `RNS_PRIME_BITS'd1116816771, `RNS_PRIME_BITS'd1998792858, `RNS_PRIME_BITS'd522676922},
    '{`RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd1022064446, `RNS_PRIME_BITS'd643203401, `RNS_PRIME_BITS'd1893865721, `RNS_PRIME_BITS'd1719835357, `RNS_PRIME_BITS'd1249075051, `RNS_PRIME_BITS'd127195022, `RNS_PRIME_BITS'd642860313, `RNS_PRIME_BITS'd1025761684, `RNS_PRIME_BITS'd2132901097, `RNS_PRIME_BITS'd320373698},
    '{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd254214852, `RNS_PRIME_BITS'd1056112510, `RNS_PRIME_BITS'd1735658448, `RNS_PRIME_BITS'd408080019, `RNS_PRIME_BITS'd886885442, `RNS_PRIME_BITS'd1702554385, `RNS_PRIME_BITS'd1984463583, `RNS_PRIME_BITS'd1228639026, `RNS_PRIME_BITS'd746257255, `RNS_PRIME_BITS'd1847365274},
    '{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1301117692, `RNS_PRIME_BITS'd121712876, `RNS_PRIME_BITS'd1725832022, `RNS_PRIME_BITS'd182045370, `RNS_PRIME_BITS'd677197750, `RNS_PRIME_BITS'd1834885785, `RNS_PRIME_BITS'd736178203, `RNS_PRIME_BITS'd507286293, `RNS_PRIME_BITS'd1266704200, `RNS_PRIME_BITS'd347681037},
    '{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd1833562202, `RNS_PRIME_BITS'd1086361181, `RNS_PRIME_BITS'd1900233247, `RNS_PRIME_BITS'd1969424525, `RNS_PRIME_BITS'd820209434, `RNS_PRIME_BITS'd324434035, `RNS_PRIME_BITS'd885531927, `RNS_PRIME_BITS'd2124779182, `RNS_PRIME_BITS'd1516624622, `RNS_PRIME_BITS'd1552400984},
    '{`RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd584132787, `RNS_PRIME_BITS'd695697577, `RNS_PRIME_BITS'd1336070358, `RNS_PRIME_BITS'd1651817411, `RNS_PRIME_BITS'd77353864, `RNS_PRIME_BITS'd1664074539, `RNS_PRIME_BITS'd1930216720, `RNS_PRIME_BITS'd1548313253, `RNS_PRIME_BITS'd598651617, `RNS_PRIME_BITS'd596604367},
    '{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd875293636, `RNS_PRIME_BITS'd2051130920, `RNS_PRIME_BITS'd421997206, `RNS_PRIME_BITS'd2060370494, `RNS_PRIME_BITS'd2144628227, `RNS_PRIME_BITS'd1566829726, `RNS_PRIME_BITS'd1386165247, `RNS_PRIME_BITS'd687714506, `RNS_PRIME_BITS'd528442972, `RNS_PRIME_BITS'd881136268},
    '{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd17774605, `RNS_PRIME_BITS'd344670759, `RNS_PRIME_BITS'd536750487, `RNS_PRIME_BITS'd221153168, `RNS_PRIME_BITS'd1979149204, `RNS_PRIME_BITS'd406483085, `RNS_PRIME_BITS'd186575011, `RNS_PRIME_BITS'd535501893, `RNS_PRIME_BITS'd1594845347, `RNS_PRIME_BITS'd724110489},
    '{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd356785962, `RNS_PRIME_BITS'd848493897, `RNS_PRIME_BITS'd1178611434, `RNS_PRIME_BITS'd905189292, `RNS_PRIME_BITS'd1769338504, `RNS_PRIME_BITS'd1348092004, `RNS_PRIME_BITS'd39071353, `RNS_PRIME_BITS'd292258251, `RNS_PRIME_BITS'd1150247224, `RNS_PRIME_BITS'd31110500},
    '{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd2038988113, `RNS_PRIME_BITS'd611046607, `RNS_PRIME_BITS'd618796859, `RNS_PRIME_BITS'd1325394714, `RNS_PRIME_BITS'd103348431, `RNS_PRIME_BITS'd997317807, `RNS_PRIME_BITS'd1569538712, `RNS_PRIME_BITS'd14021605, `RNS_PRIME_BITS'd1878121717, `RNS_PRIME_BITS'd1100880140},
    '{`RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd955160690, `RNS_PRIME_BITS'd2011563958, `RNS_PRIME_BITS'd1472788446, `RNS_PRIME_BITS'd62717420, `RNS_PRIME_BITS'd2012260124, `RNS_PRIME_BITS'd559001618, `RNS_PRIME_BITS'd1164897979, `RNS_PRIME_BITS'd999372216, `RNS_PRIME_BITS'd447044912, `RNS_PRIME_BITS'd1725572759},
    '{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd1328378368, `RNS_PRIME_BITS'd1065701949, `RNS_PRIME_BITS'd2121645181, `RNS_PRIME_BITS'd188295079, `RNS_PRIME_BITS'd2031844080, `RNS_PRIME_BITS'd1427848259, `RNS_PRIME_BITS'd1742646525, `RNS_PRIME_BITS'd1958000551, `RNS_PRIME_BITS'd690876606, `RNS_PRIME_BITS'd425238815},
    '{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd1144173285, `RNS_PRIME_BITS'd335008896, `RNS_PRIME_BITS'd1491675868, `RNS_PRIME_BITS'd776025039, `RNS_PRIME_BITS'd1631724075, `RNS_PRIME_BITS'd297212828, `RNS_PRIME_BITS'd1766860546, `RNS_PRIME_BITS'd1558486882, `RNS_PRIME_BITS'd2131064174, `RNS_PRIME_BITS'd1857760093},
    '{`RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd781130222, `RNS_PRIME_BITS'd1566302183, `RNS_PRIME_BITS'd2003607145, `RNS_PRIME_BITS'd565387027, `RNS_PRIME_BITS'd1894897721, `RNS_PRIME_BITS'd227886979, `RNS_PRIME_BITS'd1814827202, `RNS_PRIME_BITS'd835285449, `RNS_PRIME_BITS'd1573859024, `RNS_PRIME_BITS'd715601790},
    '{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd268845809, `RNS_PRIME_BITS'd816075104, `RNS_PRIME_BITS'd934272159, `RNS_PRIME_BITS'd1397979561, `RNS_PRIME_BITS'd2019979570, `RNS_PRIME_BITS'd688786362, `RNS_PRIME_BITS'd454005626, `RNS_PRIME_BITS'd2074865574, `RNS_PRIME_BITS'd2135898027, `RNS_PRIME_BITS'd1172573837},
    '{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd1825799892, `RNS_PRIME_BITS'd247813306, `RNS_PRIME_BITS'd225220907, `RNS_PRIME_BITS'd1664933581, `RNS_PRIME_BITS'd2084276684, `RNS_PRIME_BITS'd1661051490, `RNS_PRIME_BITS'd1438525080, `RNS_PRIME_BITS'd2058814547, `RNS_PRIME_BITS'd1894573574, `RNS_PRIME_BITS'd687762618},
    '{`RNS_PRIME_BITS'd213, `RNS_PRIME_BITS'd1240852021, `RNS_PRIME_BITS'd1799236445, `RNS_PRIME_BITS'd480194134, `RNS_PRIME_BITS'd448680268, `RNS_PRIME_BITS'd28101663, `RNS_PRIME_BITS'd1068560887, `RNS_PRIME_BITS'd759328019, `RNS_PRIME_BITS'd162015902, `RNS_PRIME_BITS'd1871400993, `RNS_PRIME_BITS'd1472190862},
    '{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd1464300718, `RNS_PRIME_BITS'd158825453, `RNS_PRIME_BITS'd48193229, `RNS_PRIME_BITS'd1622276664, `RNS_PRIME_BITS'd2071146701, `RNS_PRIME_BITS'd136974249, `RNS_PRIME_BITS'd1770253112, `RNS_PRIME_BITS'd1653112125, `RNS_PRIME_BITS'd1133412400, `RNS_PRIME_BITS'd69150429},
    '{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd386689036, `RNS_PRIME_BITS'd1972921725, `RNS_PRIME_BITS'd1751633961, `RNS_PRIME_BITS'd327342002, `RNS_PRIME_BITS'd1726513724, `RNS_PRIME_BITS'd857604895, `RNS_PRIME_BITS'd196079291, `RNS_PRIME_BITS'd113413555, `RNS_PRIME_BITS'd179293895, `RNS_PRIME_BITS'd100085132},
    '{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd1486183251, `RNS_PRIME_BITS'd692318239, `RNS_PRIME_BITS'd1708385398, `RNS_PRIME_BITS'd540905663, `RNS_PRIME_BITS'd568261748, `RNS_PRIME_BITS'd870281389, `RNS_PRIME_BITS'd941938269, `RNS_PRIME_BITS'd859481359, `RNS_PRIME_BITS'd1172009225, `RNS_PRIME_BITS'd614244743},
    '{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1368379953, `RNS_PRIME_BITS'd281004805, `RNS_PRIME_BITS'd29758940, `RNS_PRIME_BITS'd1956354845, `RNS_PRIME_BITS'd121223137, `RNS_PRIME_BITS'd330800609, `RNS_PRIME_BITS'd269352175, `RNS_PRIME_BITS'd1554117857, `RNS_PRIME_BITS'd438507820, `RNS_PRIME_BITS'd1830179921},
    '{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd1119124109, `RNS_PRIME_BITS'd141147247, `RNS_PRIME_BITS'd1977645907, `RNS_PRIME_BITS'd1278113227, `RNS_PRIME_BITS'd629363282, `RNS_PRIME_BITS'd2108265757, `RNS_PRIME_BITS'd332690711, `RNS_PRIME_BITS'd867978566, `RNS_PRIME_BITS'd977828196, `RNS_PRIME_BITS'd1403519540},
    '{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd1748752439, `RNS_PRIME_BITS'd581229285, `RNS_PRIME_BITS'd756157563, `RNS_PRIME_BITS'd1492554435, `RNS_PRIME_BITS'd1526862685, `RNS_PRIME_BITS'd812704507, `RNS_PRIME_BITS'd1689317871, `RNS_PRIME_BITS'd1098060407, `RNS_PRIME_BITS'd149598561, `RNS_PRIME_BITS'd1576410714},
    '{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd957539307, `RNS_PRIME_BITS'd1386640185, `RNS_PRIME_BITS'd264416368, `RNS_PRIME_BITS'd1653862382, `RNS_PRIME_BITS'd168310539, `RNS_PRIME_BITS'd980834125, `RNS_PRIME_BITS'd1648751739, `RNS_PRIME_BITS'd683132183, `RNS_PRIME_BITS'd1848768626, `RNS_PRIME_BITS'd1932282581},
    '{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1125311264, `RNS_PRIME_BITS'd389570102, `RNS_PRIME_BITS'd830221424, `RNS_PRIME_BITS'd1469660074, `RNS_PRIME_BITS'd1490586358, `RNS_PRIME_BITS'd1304060276, `RNS_PRIME_BITS'd1705708466, `RNS_PRIME_BITS'd1693472326, `RNS_PRIME_BITS'd332165351, `RNS_PRIME_BITS'd1206867073},
    '{`RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd2055724711, `RNS_PRIME_BITS'd1152721697, `RNS_PRIME_BITS'd1920620573, `RNS_PRIME_BITS'd494936011, `RNS_PRIME_BITS'd1402258395, `RNS_PRIME_BITS'd36871064, `RNS_PRIME_BITS'd1597511254, `RNS_PRIME_BITS'd1380931880, `RNS_PRIME_BITS'd1387035859, `RNS_PRIME_BITS'd746314798},
    '{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1973052422, `RNS_PRIME_BITS'd2050935508, `RNS_PRIME_BITS'd1199928760, `RNS_PRIME_BITS'd574985373, `RNS_PRIME_BITS'd1853517361, `RNS_PRIME_BITS'd1874029180, `RNS_PRIME_BITS'd1655790123, `RNS_PRIME_BITS'd225482241, `RNS_PRIME_BITS'd673834071, `RNS_PRIME_BITS'd1635235279},
    '{`RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd626565169, `RNS_PRIME_BITS'd678148867, `RNS_PRIME_BITS'd1413085432, `RNS_PRIME_BITS'd229789241, `RNS_PRIME_BITS'd669175024, `RNS_PRIME_BITS'd507705345, `RNS_PRIME_BITS'd815852633, `RNS_PRIME_BITS'd1076325068, `RNS_PRIME_BITS'd113939354, `RNS_PRIME_BITS'd1225771145},
    '{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd713461989, `RNS_PRIME_BITS'd2071007759, `RNS_PRIME_BITS'd1074126258, `RNS_PRIME_BITS'd895565421, `RNS_PRIME_BITS'd331930671, `RNS_PRIME_BITS'd540759405, `RNS_PRIME_BITS'd1934373040, `RNS_PRIME_BITS'd957049445, `RNS_PRIME_BITS'd1289346430, `RNS_PRIME_BITS'd130726263},
    '{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd33303951, `RNS_PRIME_BITS'd251669112, `RNS_PRIME_BITS'd871527458, `RNS_PRIME_BITS'd2063459396, `RNS_PRIME_BITS'd1880160642, `RNS_PRIME_BITS'd135799669, `RNS_PRIME_BITS'd1473417439, `RNS_PRIME_BITS'd1445942374, `RNS_PRIME_BITS'd858408430, `RNS_PRIME_BITS'd372366983},
    '{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd350105513, `RNS_PRIME_BITS'd961135379, `RNS_PRIME_BITS'd1546300093, `RNS_PRIME_BITS'd620076777, `RNS_PRIME_BITS'd1908843730, `RNS_PRIME_BITS'd473647087, `RNS_PRIME_BITS'd345078151, `RNS_PRIME_BITS'd1267134975, `RNS_PRIME_BITS'd1254654714, `RNS_PRIME_BITS'd1064539738},
    '{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd1455447908, `RNS_PRIME_BITS'd1972902860, `RNS_PRIME_BITS'd718563074, `RNS_PRIME_BITS'd204067039, `RNS_PRIME_BITS'd349407258, `RNS_PRIME_BITS'd2000831818, `RNS_PRIME_BITS'd74680898, `RNS_PRIME_BITS'd460758273, `RNS_PRIME_BITS'd540756407, `RNS_PRIME_BITS'd811256261},
    '{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1831138265, `RNS_PRIME_BITS'd1676556220, `RNS_PRIME_BITS'd2126107401, `RNS_PRIME_BITS'd588314791, `RNS_PRIME_BITS'd1672180200, `RNS_PRIME_BITS'd225922393, `RNS_PRIME_BITS'd328312322, `RNS_PRIME_BITS'd1084403058, `RNS_PRIME_BITS'd358945894, `RNS_PRIME_BITS'd1676468327},
    '{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd1405399662, `RNS_PRIME_BITS'd1009669518, `RNS_PRIME_BITS'd423807776, `RNS_PRIME_BITS'd1647295872, `RNS_PRIME_BITS'd1289297062, `RNS_PRIME_BITS'd856865827, `RNS_PRIME_BITS'd1387044625, `RNS_PRIME_BITS'd545736177, `RNS_PRIME_BITS'd216082995, `RNS_PRIME_BITS'd1681719117},
    '{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd184742794, `RNS_PRIME_BITS'd336386816, `RNS_PRIME_BITS'd633795346, `RNS_PRIME_BITS'd705383058, `RNS_PRIME_BITS'd1442682816, `RNS_PRIME_BITS'd412772601, `RNS_PRIME_BITS'd918401803, `RNS_PRIME_BITS'd683646684, `RNS_PRIME_BITS'd2141610068, `RNS_PRIME_BITS'd899635798},
    '{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1044496195, `RNS_PRIME_BITS'd151883032, `RNS_PRIME_BITS'd90794750, `RNS_PRIME_BITS'd731884915, `RNS_PRIME_BITS'd1867560061, `RNS_PRIME_BITS'd951019813, `RNS_PRIME_BITS'd1579805212, `RNS_PRIME_BITS'd1917741180, `RNS_PRIME_BITS'd540905734, `RNS_PRIME_BITS'd2065330097},
    '{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd761311156, `RNS_PRIME_BITS'd774727052, `RNS_PRIME_BITS'd1195992423, `RNS_PRIME_BITS'd2091990130, `RNS_PRIME_BITS'd966823518, `RNS_PRIME_BITS'd989808184, `RNS_PRIME_BITS'd1587752627, `RNS_PRIME_BITS'd1719837955, `RNS_PRIME_BITS'd1280694591, `RNS_PRIME_BITS'd662979577},
    '{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd1053061321, `RNS_PRIME_BITS'd1242808425, `RNS_PRIME_BITS'd1686683653, `RNS_PRIME_BITS'd1128449189, `RNS_PRIME_BITS'd829483264, `RNS_PRIME_BITS'd2122107396, `RNS_PRIME_BITS'd900455084, `RNS_PRIME_BITS'd933692158, `RNS_PRIME_BITS'd1329685250, `RNS_PRIME_BITS'd1050632062},
    '{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd1242777573, `RNS_PRIME_BITS'd1480771520, `RNS_PRIME_BITS'd655871583, `RNS_PRIME_BITS'd468131553, `RNS_PRIME_BITS'd1715109801, `RNS_PRIME_BITS'd1436464703, `RNS_PRIME_BITS'd1005841047, `RNS_PRIME_BITS'd356254265, `RNS_PRIME_BITS'd952212611, `RNS_PRIME_BITS'd794435263},
    '{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd519640201, `RNS_PRIME_BITS'd944885152, `RNS_PRIME_BITS'd970106672, `RNS_PRIME_BITS'd241316645, `RNS_PRIME_BITS'd1372606738, `RNS_PRIME_BITS'd2059104145, `RNS_PRIME_BITS'd679179388, `RNS_PRIME_BITS'd1492041218, `RNS_PRIME_BITS'd1824216637, `RNS_PRIME_BITS'd66648376},
    '{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd1978003332, `RNS_PRIME_BITS'd478263574, `RNS_PRIME_BITS'd1785392179, `RNS_PRIME_BITS'd1197953276, `RNS_PRIME_BITS'd106057337, `RNS_PRIME_BITS'd2145826994, `RNS_PRIME_BITS'd205573307, `RNS_PRIME_BITS'd947890726, `RNS_PRIME_BITS'd1094961097, `RNS_PRIME_BITS'd720404290},
    '{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd1147003102, `RNS_PRIME_BITS'd221482402, `RNS_PRIME_BITS'd1824474512, `RNS_PRIME_BITS'd519041421, `RNS_PRIME_BITS'd673860316, `RNS_PRIME_BITS'd180340212, `RNS_PRIME_BITS'd1018677988, `RNS_PRIME_BITS'd1821615501, `RNS_PRIME_BITS'd2122077440, `RNS_PRIME_BITS'd309168117},
    '{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd12870039, `RNS_PRIME_BITS'd278774359, `RNS_PRIME_BITS'd999290885, `RNS_PRIME_BITS'd1746389166, `RNS_PRIME_BITS'd206584424, `RNS_PRIME_BITS'd815127430, `RNS_PRIME_BITS'd343227041, `RNS_PRIME_BITS'd508295792, `RNS_PRIME_BITS'd451346596, `RNS_PRIME_BITS'd1604242461},
    '{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1358866390, `RNS_PRIME_BITS'd1534498320, `RNS_PRIME_BITS'd108997519, `RNS_PRIME_BITS'd1478988427, `RNS_PRIME_BITS'd2022885132, `RNS_PRIME_BITS'd1564793906, `RNS_PRIME_BITS'd1443506900, `RNS_PRIME_BITS'd1015344614, `RNS_PRIME_BITS'd617070652, `RNS_PRIME_BITS'd1829857110},
    '{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd694384824, `RNS_PRIME_BITS'd2033364169, `RNS_PRIME_BITS'd453130443, `RNS_PRIME_BITS'd1758966300, `RNS_PRIME_BITS'd974564895, `RNS_PRIME_BITS'd948406233, `RNS_PRIME_BITS'd1121340545, `RNS_PRIME_BITS'd1724578302, `RNS_PRIME_BITS'd381422488, `RNS_PRIME_BITS'd982359344},
    '{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd967763240, `RNS_PRIME_BITS'd1427971716, `RNS_PRIME_BITS'd494910485, `RNS_PRIME_BITS'd492740892, `RNS_PRIME_BITS'd273173563, `RNS_PRIME_BITS'd658460783, `RNS_PRIME_BITS'd2080148280, `RNS_PRIME_BITS'd621597327, `RNS_PRIME_BITS'd1943862185, `RNS_PRIME_BITS'd326449776},
    '{`RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd1675838128, `RNS_PRIME_BITS'd468707300, `RNS_PRIME_BITS'd799885904, `RNS_PRIME_BITS'd1854190662, `RNS_PRIME_BITS'd268681678, `RNS_PRIME_BITS'd1719671837, `RNS_PRIME_BITS'd1282259653, `RNS_PRIME_BITS'd744227196, `RNS_PRIME_BITS'd3314132, `RNS_PRIME_BITS'd1601120085},
    '{`RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd1614885743, `RNS_PRIME_BITS'd1859106025, `RNS_PRIME_BITS'd625570152, `RNS_PRIME_BITS'd866216548, `RNS_PRIME_BITS'd1641084080, `RNS_PRIME_BITS'd737429472, `RNS_PRIME_BITS'd1677505507, `RNS_PRIME_BITS'd735874166, `RNS_PRIME_BITS'd712493476, `RNS_PRIME_BITS'd475235749},
    '{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd577663718, `RNS_PRIME_BITS'd1235052902, `RNS_PRIME_BITS'd1798892458, `RNS_PRIME_BITS'd1499030155, `RNS_PRIME_BITS'd1774223663, `RNS_PRIME_BITS'd1714899668, `RNS_PRIME_BITS'd1902694704, `RNS_PRIME_BITS'd936281940, `RNS_PRIME_BITS'd670751538, `RNS_PRIME_BITS'd97394646},
    '{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1655002074, `RNS_PRIME_BITS'd1377669667, `RNS_PRIME_BITS'd1984677102, `RNS_PRIME_BITS'd1793490330, `RNS_PRIME_BITS'd355605847, `RNS_PRIME_BITS'd1512149371, `RNS_PRIME_BITS'd1564130907, `RNS_PRIME_BITS'd1144315676, `RNS_PRIME_BITS'd593371229, `RNS_PRIME_BITS'd991236607}
};

parameter B_BASIS_poly twist_factor_b   = '{
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1},
    '{`RNS_PRIME_BITS'd982714381, `RNS_PRIME_BITS'd561201457, `RNS_PRIME_BITS'd2030504833, `RNS_PRIME_BITS'd520071954, `RNS_PRIME_BITS'd1910348564, `RNS_PRIME_BITS'd1111366840, `RNS_PRIME_BITS'd1316470784, `RNS_PRIME_BITS'd2130228297, `RNS_PRIME_BITS'd1972786723, `RNS_PRIME_BITS'd601347331},
    '{`RNS_PRIME_BITS'd1654849230, `RNS_PRIME_BITS'd318222520, `RNS_PRIME_BITS'd458644985, `RNS_PRIME_BITS'd1659477478, `RNS_PRIME_BITS'd221897449, `RNS_PRIME_BITS'd1817702166, `RNS_PRIME_BITS'd1453892451, `RNS_PRIME_BITS'd1033346514, `RNS_PRIME_BITS'd1445995283, `RNS_PRIME_BITS'd330138710},
    '{`RNS_PRIME_BITS'd478051828, `RNS_PRIME_BITS'd1438809348, `RNS_PRIME_BITS'd1933006424, `RNS_PRIME_BITS'd380013956, `RNS_PRIME_BITS'd367995126, `RNS_PRIME_BITS'd308654393, `RNS_PRIME_BITS'd1313726466, `RNS_PRIME_BITS'd581750232, `RNS_PRIME_BITS'd1987253116, `RNS_PRIME_BITS'd1006948292},
    '{`RNS_PRIME_BITS'd356657619, `RNS_PRIME_BITS'd1828267041, `RNS_PRIME_BITS'd2042051371, `RNS_PRIME_BITS'd532048860, `RNS_PRIME_BITS'd1539132485, `RNS_PRIME_BITS'd1902036916, `RNS_PRIME_BITS'd1435226373, `RNS_PRIME_BITS'd1625142860, `RNS_PRIME_BITS'd501746762, `RNS_PRIME_BITS'd211376156},
    '{`RNS_PRIME_BITS'd1920663579, `RNS_PRIME_BITS'd1617885585, `RNS_PRIME_BITS'd734171544, `RNS_PRIME_BITS'd1587022193, `RNS_PRIME_BITS'd2051390243, `RNS_PRIME_BITS'd1514881435, `RNS_PRIME_BITS'd789663591, `RNS_PRIME_BITS'd486721859, `RNS_PRIME_BITS'd463114787, `RNS_PRIME_BITS'd15801270},
    '{`RNS_PRIME_BITS'd302866737, `RNS_PRIME_BITS'd1310190713, `RNS_PRIME_BITS'd2001209167, `RNS_PRIME_BITS'd678117384, `RNS_PRIME_BITS'd2024510820, `RNS_PRIME_BITS'd203341575, `RNS_PRIME_BITS'd1428696568, `RNS_PRIME_BITS'd571204460, `RNS_PRIME_BITS'd108107719, `RNS_PRIME_BITS'd97888807},
    '{`RNS_PRIME_BITS'd351262005, `RNS_PRIME_BITS'd1915188815, `RNS_PRIME_BITS'd1270889040, `RNS_PRIME_BITS'd646964512, `RNS_PRIME_BITS'd1441807459, `RNS_PRIME_BITS'd1364034874, `RNS_PRIME_BITS'd1692753891, `RNS_PRIME_BITS'd981144746, `RNS_PRIME_BITS'd1680185572, `RNS_PRIME_BITS'd1297233476},
    '{`RNS_PRIME_BITS'd532016628, `RNS_PRIME_BITS'd1346436954, `RNS_PRIME_BITS'd662532888, `RNS_PRIME_BITS'd1599846131, `RNS_PRIME_BITS'd2041325775, `RNS_PRIME_BITS'd1781417128, `RNS_PRIME_BITS'd1222739369, `RNS_PRIME_BITS'd574229214, `RNS_PRIME_BITS'd1267807369, `RNS_PRIME_BITS'd125361803},
    '{`RNS_PRIME_BITS'd1151501468, `RNS_PRIME_BITS'd804641710, `RNS_PRIME_BITS'd332110078, `RNS_PRIME_BITS'd492774328, `RNS_PRIME_BITS'd101596083, `RNS_PRIME_BITS'd1866997580, `RNS_PRIME_BITS'd1601511596, `RNS_PRIME_BITS'd1089218493, `RNS_PRIME_BITS'd1018407763, `RNS_PRIME_BITS'd1327782020},
    '{`RNS_PRIME_BITS'd652946039, `RNS_PRIME_BITS'd1430678598, `RNS_PRIME_BITS'd586122886, `RNS_PRIME_BITS'd1813223460, `RNS_PRIME_BITS'd411860025, `RNS_PRIME_BITS'd337893308, `RNS_PRIME_BITS'd1424810859, `RNS_PRIME_BITS'd26513139, `RNS_PRIME_BITS'd1846795101, `RNS_PRIME_BITS'd774401595},
    '{`RNS_PRIME_BITS'd1144091943, `RNS_PRIME_BITS'd1654629824, `RNS_PRIME_BITS'd1868204885, `RNS_PRIME_BITS'd2035977623, `RNS_PRIME_BITS'd1825753344, `RNS_PRIME_BITS'd859229142, `RNS_PRIME_BITS'd1150701755, `RNS_PRIME_BITS'd2010605865, `RNS_PRIME_BITS'd1267530456, `RNS_PRIME_BITS'd993630259},
    '{`RNS_PRIME_BITS'd1233595480, `RNS_PRIME_BITS'd400618345, `RNS_PRIME_BITS'd633289293, `RNS_PRIME_BITS'd451198491, `RNS_PRIME_BITS'd1284434959, `RNS_PRIME_BITS'd181333865, `RNS_PRIME_BITS'd1443308359, `RNS_PRIME_BITS'd341692242, `RNS_PRIME_BITS'd246731728, `RNS_PRIME_BITS'd830621476},
    '{`RNS_PRIME_BITS'd327413943, `RNS_PRIME_BITS'd1866406664, `RNS_PRIME_BITS'd1828476394, `RNS_PRIME_BITS'd1649721566, `RNS_PRIME_BITS'd341435820, `RNS_PRIME_BITS'd162479211, `RNS_PRIME_BITS'd214516484, `RNS_PRIME_BITS'd1506386962, `RNS_PRIME_BITS'd1125681298, `RNS_PRIME_BITS'd213719977},
    '{`RNS_PRIME_BITS'd849304041, `RNS_PRIME_BITS'd5588299, `RNS_PRIME_BITS'd1282347525, `RNS_PRIME_BITS'd2112063758, `RNS_PRIME_BITS'd323800841, `RNS_PRIME_BITS'd1144062347, `RNS_PRIME_BITS'd908740576, `RNS_PRIME_BITS'd1816898220, `RNS_PRIME_BITS'd1797675798, `RNS_PRIME_BITS'd1784673181},
    '{`RNS_PRIME_BITS'd385268797, `RNS_PRIME_BITS'd120346045, `RNS_PRIME_BITS'd679192186, `RNS_PRIME_BITS'd730453618, `RNS_PRIME_BITS'd959857878, `RNS_PRIME_BITS'd1296633865, `RNS_PRIME_BITS'd918632540, `RNS_PRIME_BITS'd313660301, `RNS_PRIME_BITS'd1117135201, `RNS_PRIME_BITS'd244734214},
    '{`RNS_PRIME_BITS'd1929740512, `RNS_PRIME_BITS'd80763692, `RNS_PRIME_BITS'd1110746654, `RNS_PRIME_BITS'd1888511225, `RNS_PRIME_BITS'd747078255, `RNS_PRIME_BITS'd1071833897, `RNS_PRIME_BITS'd1181774526, `RNS_PRIME_BITS'd1944313893, `RNS_PRIME_BITS'd849564324, `RNS_PRIME_BITS'd634071871},
    '{`RNS_PRIME_BITS'd1437307346, `RNS_PRIME_BITS'd545997482, `RNS_PRIME_BITS'd1048891790, `RNS_PRIME_BITS'd1946521804, `RNS_PRIME_BITS'd172892730, `RNS_PRIME_BITS'd1132496960, `RNS_PRIME_BITS'd95042921, `RNS_PRIME_BITS'd1484566497, `RNS_PRIME_BITS'd1508207091, `RNS_PRIME_BITS'd1357050316},
    '{`RNS_PRIME_BITS'd1054516963, `RNS_PRIME_BITS'd983104082, `RNS_PRIME_BITS'd595179583, `RNS_PRIME_BITS'd1078093079, `RNS_PRIME_BITS'd1581201429, `RNS_PRIME_BITS'd265094956, `RNS_PRIME_BITS'd162700068, `RNS_PRIME_BITS'd1541045115, `RNS_PRIME_BITS'd251058699, `RNS_PRIME_BITS'd850930788},
    '{`RNS_PRIME_BITS'd2052121271, `RNS_PRIME_BITS'd2097368234, `RNS_PRIME_BITS'd1124820764, `RNS_PRIME_BITS'd1326701425, `RNS_PRIME_BITS'd285618846, `RNS_PRIME_BITS'd1422611, `RNS_PRIME_BITS'd922037797, `RNS_PRIME_BITS'd630923484, `RNS_PRIME_BITS'd1729285507, `RNS_PRIME_BITS'd1908735073},
    '{`RNS_PRIME_BITS'd470080841, `RNS_PRIME_BITS'd918812250, `RNS_PRIME_BITS'd1315499404, `RNS_PRIME_BITS'd734192161, `RNS_PRIME_BITS'd498026890, `RNS_PRIME_BITS'd536379334, `RNS_PRIME_BITS'd608940391, `RNS_PRIME_BITS'd2064395269, `RNS_PRIME_BITS'd796429192, `RNS_PRIME_BITS'd855303704},
    '{`RNS_PRIME_BITS'd1579045017, `RNS_PRIME_BITS'd2055579709, `RNS_PRIME_BITS'd674452159, `RNS_PRIME_BITS'd1770001053, `RNS_PRIME_BITS'd1516662357, `RNS_PRIME_BITS'd1941747448, `RNS_PRIME_BITS'd1162784154, `RNS_PRIME_BITS'd1090276043, `RNS_PRIME_BITS'd2067686905, `RNS_PRIME_BITS'd892337725},
    '{`RNS_PRIME_BITS'd297821259, `RNS_PRIME_BITS'd1980041940, `RNS_PRIME_BITS'd1801404655, `RNS_PRIME_BITS'd1913561989, `RNS_PRIME_BITS'd743336322, `RNS_PRIME_BITS'd987777415, `RNS_PRIME_BITS'd385218143, `RNS_PRIME_BITS'd2012553244, `RNS_PRIME_BITS'd1979833503, `RNS_PRIME_BITS'd518922129},
    '{`RNS_PRIME_BITS'd641843845, `RNS_PRIME_BITS'd1139003082, `RNS_PRIME_BITS'd1493917469, `RNS_PRIME_BITS'd965099418, `RNS_PRIME_BITS'd221590400, `RNS_PRIME_BITS'd1196073590, `RNS_PRIME_BITS'd789327398, `RNS_PRIME_BITS'd1510469846, `RNS_PRIME_BITS'd270694143, `RNS_PRIME_BITS'd120244624},
    '{`RNS_PRIME_BITS'd99841913, `RNS_PRIME_BITS'd159606694, `RNS_PRIME_BITS'd1314416481, `RNS_PRIME_BITS'd2125349561, `RNS_PRIME_BITS'd807294136, `RNS_PRIME_BITS'd2062390131, `RNS_PRIME_BITS'd1394307591, `RNS_PRIME_BITS'd337677835, `RNS_PRIME_BITS'd132886023, `RNS_PRIME_BITS'd590119148},
    '{`RNS_PRIME_BITS'd444118214, `RNS_PRIME_BITS'd820749293, `RNS_PRIME_BITS'd1952643917, `RNS_PRIME_BITS'd2020087064, `RNS_PRIME_BITS'd1720419235, `RNS_PRIME_BITS'd1850634582, `RNS_PRIME_BITS'd541471192, `RNS_PRIME_BITS'd1602631169, `RNS_PRIME_BITS'd1160547813, `RNS_PRIME_BITS'd1858954969},
    '{`RNS_PRIME_BITS'd1094401579, `RNS_PRIME_BITS'd1979993210, `RNS_PRIME_BITS'd1368761486, `RNS_PRIME_BITS'd1790284840, `RNS_PRIME_BITS'd2108289477, `RNS_PRIME_BITS'd1033810328, `RNS_PRIME_BITS'd385488776, `RNS_PRIME_BITS'd972301580, `RNS_PRIME_BITS'd464279201, `RNS_PRIME_BITS'd627138487},
    '{`RNS_PRIME_BITS'd936096522, `RNS_PRIME_BITS'd2126679887, `RNS_PRIME_BITS'd190758143, `RNS_PRIME_BITS'd653091537, `RNS_PRIME_BITS'd1402153400, `RNS_PRIME_BITS'd1801237427, `RNS_PRIME_BITS'd871114005, `RNS_PRIME_BITS'd1727682728, `RNS_PRIME_BITS'd1152260240, `RNS_PRIME_BITS'd886133038},
    '{`RNS_PRIME_BITS'd123364587, `RNS_PRIME_BITS'd229579563, `RNS_PRIME_BITS'd1292695071, `RNS_PRIME_BITS'd131782201, `RNS_PRIME_BITS'd1557026756, `RNS_PRIME_BITS'd1520994666, `RNS_PRIME_BITS'd1975029035, `RNS_PRIME_BITS'd1168805901, `RNS_PRIME_BITS'd422202768, `RNS_PRIME_BITS'd44695371},
    '{`RNS_PRIME_BITS'd456798682, `RNS_PRIME_BITS'd1169203214, `RNS_PRIME_BITS'd326439411, `RNS_PRIME_BITS'd1893247609, `RNS_PRIME_BITS'd486052227, `RNS_PRIME_BITS'd1746039191, `RNS_PRIME_BITS'd953927283, `RNS_PRIME_BITS'd1956709734, `RNS_PRIME_BITS'd48756347, `RNS_PRIME_BITS'd747272326},
    '{`RNS_PRIME_BITS'd371148888, `RNS_PRIME_BITS'd1458564334, `RNS_PRIME_BITS'd517075660, `RNS_PRIME_BITS'd303751980, `RNS_PRIME_BITS'd639432542, `RNS_PRIME_BITS'd729791605, `RNS_PRIME_BITS'd220568782, `RNS_PRIME_BITS'd73418631, `RNS_PRIME_BITS'd1842850055, `RNS_PRIME_BITS'd1029685765},
    '{`RNS_PRIME_BITS'd958225700, `RNS_PRIME_BITS'd1357775805, `RNS_PRIME_BITS'd611103098, `RNS_PRIME_BITS'd1334847884, `RNS_PRIME_BITS'd566734447, `RNS_PRIME_BITS'd1779837071, `RNS_PRIME_BITS'd1814090713, `RNS_PRIME_BITS'd1880750118, `RNS_PRIME_BITS'd583666609, `RNS_PRIME_BITS'd1598964437},
    '{`RNS_PRIME_BITS'd368900981, `RNS_PRIME_BITS'd1776948932, `RNS_PRIME_BITS'd584149928, `RNS_PRIME_BITS'd873118585, `RNS_PRIME_BITS'd1361170515, `RNS_PRIME_BITS'd1162711167, `RNS_PRIME_BITS'd2018759315, `RNS_PRIME_BITS'd2098452362, `RNS_PRIME_BITS'd1282120144, `RNS_PRIME_BITS'd764279395},
    '{`RNS_PRIME_BITS'd906812118, `RNS_PRIME_BITS'd1955170315, `RNS_PRIME_BITS'd140317819, `RNS_PRIME_BITS'd249386706, `RNS_PRIME_BITS'd1756055478, `RNS_PRIME_BITS'd915333332, `RNS_PRIME_BITS'd1392338561, `RNS_PRIME_BITS'd554672634, `RNS_PRIME_BITS'd1803248469, `RNS_PRIME_BITS'd973858991},
    '{`RNS_PRIME_BITS'd27942223, `RNS_PRIME_BITS'd1966586531, `RNS_PRIME_BITS'd855293400, `RNS_PRIME_BITS'd2042384205, `RNS_PRIME_BITS'd1707467875, `RNS_PRIME_BITS'd1299152479, `RNS_PRIME_BITS'd1860847603, `RNS_PRIME_BITS'd1726140753, `RNS_PRIME_BITS'd327226555, `RNS_PRIME_BITS'd1314367513},
    '{`RNS_PRIME_BITS'd895294767, `RNS_PRIME_BITS'd110672867, `RNS_PRIME_BITS'd714603448, `RNS_PRIME_BITS'd1211271110, `RNS_PRIME_BITS'd1147352387, `RNS_PRIME_BITS'd1301194870, `RNS_PRIME_BITS'd987706370, `RNS_PRIME_BITS'd54660901, `RNS_PRIME_BITS'd819125480, `RNS_PRIME_BITS'd1786870076},
    '{`RNS_PRIME_BITS'd1022769805, `RNS_PRIME_BITS'd1050480888, `RNS_PRIME_BITS'd1486683312, `RNS_PRIME_BITS'd499906752, `RNS_PRIME_BITS'd1986920445, `RNS_PRIME_BITS'd1980475697, `RNS_PRIME_BITS'd587044175, `RNS_PRIME_BITS'd818416481, `RNS_PRIME_BITS'd35025808, `RNS_PRIME_BITS'd996800473},
    '{`RNS_PRIME_BITS'd1552017062, `RNS_PRIME_BITS'd1649403189, `RNS_PRIME_BITS'd240212080, `RNS_PRIME_BITS'd1757234669, `RNS_PRIME_BITS'd594637207, `RNS_PRIME_BITS'd988918344, `RNS_PRIME_BITS'd99971581, `RNS_PRIME_BITS'd1747488468, `RNS_PRIME_BITS'd1882163270, `RNS_PRIME_BITS'd456097637},
    '{`RNS_PRIME_BITS'd51446398, `RNS_PRIME_BITS'd554085691, `RNS_PRIME_BITS'd840596094, `RNS_PRIME_BITS'd393905830, `RNS_PRIME_BITS'd1120665741, `RNS_PRIME_BITS'd881125819, `RNS_PRIME_BITS'd649424080, `RNS_PRIME_BITS'd1455471245, `RNS_PRIME_BITS'd458116540, `RNS_PRIME_BITS'd1687641260},
    '{`RNS_PRIME_BITS'd199576301, `RNS_PRIME_BITS'd775123075, `RNS_PRIME_BITS'd368477724, `RNS_PRIME_BITS'd1693926536, `RNS_PRIME_BITS'd914203855, `RNS_PRIME_BITS'd237869749, `RNS_PRIME_BITS'd815239180, `RNS_PRIME_BITS'd692845039, `RNS_PRIME_BITS'd768852906, `RNS_PRIME_BITS'd460818202},
    '{`RNS_PRIME_BITS'd1898245248, `RNS_PRIME_BITS'd1464394521, `RNS_PRIME_BITS'd732592157, `RNS_PRIME_BITS'd780663828, `RNS_PRIME_BITS'd1967509349, `RNS_PRIME_BITS'd1814328256, `RNS_PRIME_BITS'd216334037, `RNS_PRIME_BITS'd551036518, `RNS_PRIME_BITS'd1945334986, `RNS_PRIME_BITS'd1264514118},
    '{`RNS_PRIME_BITS'd1467943930, `RNS_PRIME_BITS'd1992441198, `RNS_PRIME_BITS'd1047139254, `RNS_PRIME_BITS'd329767801, `RNS_PRIME_BITS'd1977879822, `RNS_PRIME_BITS'd627285491, `RNS_PRIME_BITS'd1040898177, `RNS_PRIME_BITS'd1927967098, `RNS_PRIME_BITS'd1632011555, `RNS_PRIME_BITS'd1401930789},
    '{`RNS_PRIME_BITS'd1732476368, `RNS_PRIME_BITS'd1295673068, `RNS_PRIME_BITS'd1079673294, `RNS_PRIME_BITS'd2044280699, `RNS_PRIME_BITS'd1932873997, `RNS_PRIME_BITS'd718059950, `RNS_PRIME_BITS'd1226695548, `RNS_PRIME_BITS'd319374927, `RNS_PRIME_BITS'd1006104391, `RNS_PRIME_BITS'd703232155},
    '{`RNS_PRIME_BITS'd559257721, `RNS_PRIME_BITS'd1767109925, `RNS_PRIME_BITS'd1351312793, `RNS_PRIME_BITS'd379354092, `RNS_PRIME_BITS'd902553616, `RNS_PRIME_BITS'd1567408049, `RNS_PRIME_BITS'd2004174612, `RNS_PRIME_BITS'd1915883062, `RNS_PRIME_BITS'd1568208839, `RNS_PRIME_BITS'd799915249},
    '{`RNS_PRIME_BITS'd1631487701, `RNS_PRIME_BITS'd1096154473, `RNS_PRIME_BITS'd1594888548, `RNS_PRIME_BITS'd1987906920, `RNS_PRIME_BITS'd1275904696, `RNS_PRIME_BITS'd45733247, `RNS_PRIME_BITS'd2109392002, `RNS_PRIME_BITS'd1049625500, `RNS_PRIME_BITS'd1719836841, `RNS_PRIME_BITS'd279176347},
    '{`RNS_PRIME_BITS'd1721817336, `RNS_PRIME_BITS'd767563666, `RNS_PRIME_BITS'd1273959981, `RNS_PRIME_BITS'd1075761591, `RNS_PRIME_BITS'd187303824, `RNS_PRIME_BITS'd1822384920, `RNS_PRIME_BITS'd133379464, `RNS_PRIME_BITS'd184438272, `RNS_PRIME_BITS'd1461368271, `RNS_PRIME_BITS'd313264892},
    '{`RNS_PRIME_BITS'd421878258, `RNS_PRIME_BITS'd674822329, `RNS_PRIME_BITS'd196565656, `RNS_PRIME_BITS'd1790217672, `RNS_PRIME_BITS'd1691018214, `RNS_PRIME_BITS'd1758326586, `RNS_PRIME_BITS'd1733682231, `RNS_PRIME_BITS'd1734877556, `RNS_PRIME_BITS'd416072182, `RNS_PRIME_BITS'd1441277666},
    '{`RNS_PRIME_BITS'd557994804, `RNS_PRIME_BITS'd1072848871, `RNS_PRIME_BITS'd1394641272, `RNS_PRIME_BITS'd1753588508, `RNS_PRIME_BITS'd2146447664, `RNS_PRIME_BITS'd1454548222, `RNS_PRIME_BITS'd2118490453, `RNS_PRIME_BITS'd1685711725, `RNS_PRIME_BITS'd726102973, `RNS_PRIME_BITS'd223845845},
    '{`RNS_PRIME_BITS'd304649431, `RNS_PRIME_BITS'd552851043, `RNS_PRIME_BITS'd500041537, `RNS_PRIME_BITS'd2052067642, `RNS_PRIME_BITS'd2080135103, `RNS_PRIME_BITS'd1467683836, `RNS_PRIME_BITS'd353404950, `RNS_PRIME_BITS'd1945521432, `RNS_PRIME_BITS'd1970029940, `RNS_PRIME_BITS'd2061554458},
    '{`RNS_PRIME_BITS'd8907008, `RNS_PRIME_BITS'd1274432900, `RNS_PRIME_BITS'd713754135, `RNS_PRIME_BITS'd88328166, `RNS_PRIME_BITS'd690462842, `RNS_PRIME_BITS'd630505524, `RNS_PRIME_BITS'd286276109, `RNS_PRIME_BITS'd1094799911, `RNS_PRIME_BITS'd1229835195, `RNS_PRIME_BITS'd1665960726},
    '{`RNS_PRIME_BITS'd271032415, `RNS_PRIME_BITS'd1263489667, `RNS_PRIME_BITS'd1873914868, `RNS_PRIME_BITS'd102380589, `RNS_PRIME_BITS'd466893867, `RNS_PRIME_BITS'd275250926, `RNS_PRIME_BITS'd86404339, `RNS_PRIME_BITS'd353031189, `RNS_PRIME_BITS'd611355256, `RNS_PRIME_BITS'd990739525},
    '{`RNS_PRIME_BITS'd1720040104, `RNS_PRIME_BITS'd885989717, `RNS_PRIME_BITS'd1078246245, `RNS_PRIME_BITS'd1561618962, `RNS_PRIME_BITS'd1038541210, `RNS_PRIME_BITS'd770159278, `RNS_PRIME_BITS'd1246377055, `RNS_PRIME_BITS'd1813434134, `RNS_PRIME_BITS'd792897446, `RNS_PRIME_BITS'd76817238},
    '{`RNS_PRIME_BITS'd1766152386, `RNS_PRIME_BITS'd236666624, `RNS_PRIME_BITS'd514903787, `RNS_PRIME_BITS'd1443630163, `RNS_PRIME_BITS'd1022960172, `RNS_PRIME_BITS'd1343151649, `RNS_PRIME_BITS'd972264218, `RNS_PRIME_BITS'd1923012750, `RNS_PRIME_BITS'd108303762, `RNS_PRIME_BITS'd616062626},
    '{`RNS_PRIME_BITS'd809081996, `RNS_PRIME_BITS'd1923634752, `RNS_PRIME_BITS'd1737225677, `RNS_PRIME_BITS'd1636333534, `RNS_PRIME_BITS'd1108497895, `RNS_PRIME_BITS'd136842044, `RNS_PRIME_BITS'd350723734, `RNS_PRIME_BITS'd1158896720, `RNS_PRIME_BITS'd928987687, `RNS_PRIME_BITS'd1278419481},
    '{`RNS_PRIME_BITS'd1651675396, `RNS_PRIME_BITS'd147052478, `RNS_PRIME_BITS'd1438162619, `RNS_PRIME_BITS'd2056193828, `RNS_PRIME_BITS'd171133878, `RNS_PRIME_BITS'd103088552, `RNS_PRIME_BITS'd611788180, `RNS_PRIME_BITS'd1273570555, `RNS_PRIME_BITS'd2141801975, `RNS_PRIME_BITS'd1138746994},
    '{`RNS_PRIME_BITS'd1331311885, `RNS_PRIME_BITS'd773740556, `RNS_PRIME_BITS'd1755701290, `RNS_PRIME_BITS'd1878383483, `RNS_PRIME_BITS'd1121975700, `RNS_PRIME_BITS'd898174659, `RNS_PRIME_BITS'd2046419506, `RNS_PRIME_BITS'd130023201, `RNS_PRIME_BITS'd1602925057, `RNS_PRIME_BITS'd740347681},
    '{`RNS_PRIME_BITS'd769115895, `RNS_PRIME_BITS'd1915037, `RNS_PRIME_BITS'd657916126, `RNS_PRIME_BITS'd763768649, `RNS_PRIME_BITS'd1239138918, `RNS_PRIME_BITS'd218696274, `RNS_PRIME_BITS'd211766403, `RNS_PRIME_BITS'd1362281852, `RNS_PRIME_BITS'd1719197983, `RNS_PRIME_BITS'd794875457},
    '{`RNS_PRIME_BITS'd1990768752, `RNS_PRIME_BITS'd1795377192, `RNS_PRIME_BITS'd743489674, `RNS_PRIME_BITS'd1663859725, `RNS_PRIME_BITS'd58964999, `RNS_PRIME_BITS'd1758502347, `RNS_PRIME_BITS'd1172996175, `RNS_PRIME_BITS'd96243187, `RNS_PRIME_BITS'd1842468980, `RNS_PRIME_BITS'd1779277119},
    '{`RNS_PRIME_BITS'd1644425917, `RNS_PRIME_BITS'd674188376, `RNS_PRIME_BITS'd970993592, `RNS_PRIME_BITS'd1883950119, `RNS_PRIME_BITS'd1584543981, `RNS_PRIME_BITS'd194569702, `RNS_PRIME_BITS'd1142519638, `RNS_PRIME_BITS'd1736961913, `RNS_PRIME_BITS'd335514896, `RNS_PRIME_BITS'd1006865747},
    '{`RNS_PRIME_BITS'd1206592301, `RNS_PRIME_BITS'd1038169980, `RNS_PRIME_BITS'd1544729701, `RNS_PRIME_BITS'd1765983319, `RNS_PRIME_BITS'd1014783106, `RNS_PRIME_BITS'd1833115473, `RNS_PRIME_BITS'd93701488, `RNS_PRIME_BITS'd1821585998, `RNS_PRIME_BITS'd1974242872, `RNS_PRIME_BITS'd1512458516},
    '{`RNS_PRIME_BITS'd1688834505, `RNS_PRIME_BITS'd155056032, `RNS_PRIME_BITS'd677137612, `RNS_PRIME_BITS'd1170752224, `RNS_PRIME_BITS'd319429885, `RNS_PRIME_BITS'd2146875856, `RNS_PRIME_BITS'd1943881058, `RNS_PRIME_BITS'd695913565, `RNS_PRIME_BITS'd1405654688, `RNS_PRIME_BITS'd520640850},
    '{`RNS_PRIME_BITS'd1022667949, `RNS_PRIME_BITS'd1063723561, `RNS_PRIME_BITS'd1980951143, `RNS_PRIME_BITS'd1028658040, `RNS_PRIME_BITS'd77300856, `RNS_PRIME_BITS'd1385487051, `RNS_PRIME_BITS'd1817397096, `RNS_PRIME_BITS'd694079929, `RNS_PRIME_BITS'd1947249161, `RNS_PRIME_BITS'd629079252},
    '{`RNS_PRIME_BITS'd826531416, `RNS_PRIME_BITS'd552348229, `RNS_PRIME_BITS'd1474472800, `RNS_PRIME_BITS'd581664342, `RNS_PRIME_BITS'd2100968896, `RNS_PRIME_BITS'd594047528, `RNS_PRIME_BITS'd752878080, `RNS_PRIME_BITS'd295372288, `RNS_PRIME_BITS'd862305235, `RNS_PRIME_BITS'd1708924581},
    '{`RNS_PRIME_BITS'd423155928, `RNS_PRIME_BITS'd2022047502, `RNS_PRIME_BITS'd895771398, `RNS_PRIME_BITS'd164737598, `RNS_PRIME_BITS'd538728578, `RNS_PRIME_BITS'd91096341, `RNS_PRIME_BITS'd1545542847, `RNS_PRIME_BITS'd592953865, `RNS_PRIME_BITS'd516818747, `RNS_PRIME_BITS'd1490950549}
};
parameter B_BASIS_poly untwist_factor_b =  '{
    '{`RNS_PRIME_BITS'd2113938037, `RNS_PRIME_BITS'd2113939297, `RNS_PRIME_BITS'd2113939675, `RNS_PRIME_BITS'd2113939927, `RNS_PRIME_BITS'd2113940305, `RNS_PRIME_BITS'd2113941061, `RNS_PRIME_BITS'd2113941565, `RNS_PRIME_BITS'd2113942321, `RNS_PRIME_BITS'd2113944841, `RNS_PRIME_BITS'd2113947613},
    '{`RNS_PRIME_BITS'd798697917, `RNS_PRIME_BITS'd438169796, `RNS_PRIME_BITS'd187331160, `RNS_PRIME_BITS'd2077811300, `RNS_PRIME_BITS'd58691582, `RNS_PRIME_BITS'd703223640, `RNS_PRIME_BITS'd2089792458, `RNS_PRIME_BITS'd292726856, `RNS_PRIME_BITS'd1971650828, `RNS_PRIME_BITS'd681353102},
    '{`RNS_PRIME_BITS'd792395175, `RNS_PRIME_BITS'd159142519, `RNS_PRIME_BITS'd1050708499, `RNS_PRIME_BITS'd729112739, `RNS_PRIME_BITS'd2114667274, `RNS_PRIME_BITS'd1332902808, `RNS_PRIME_BITS'd2135732473, `RNS_PRIME_BITS'd2142881769, `RNS_PRIME_BITS'd624065401, `RNS_PRIME_BITS'd1214822842},
    '{`RNS_PRIME_BITS'd1493976554, `RNS_PRIME_BITS'd1359117592, `RNS_PRIME_BITS'd1277676961, `RNS_PRIME_BITS'd1862984931, `RNS_PRIME_BITS'd1877850223, `RNS_PRIME_BITS'd347452585, `RNS_PRIME_BITS'd1313788291, `RNS_PRIME_BITS'd1901769482, `RNS_PRIME_BITS'd271566352, `RNS_PRIME_BITS'd661265117},
    '{`RNS_PRIME_BITS'd275603109, `RNS_PRIME_BITS'd1071324194, `RNS_PRIME_BITS'd392074901, `RNS_PRIME_BITS'd1055454261, `RNS_PRIME_BITS'd2041839997, `RNS_PRIME_BITS'd503328985, `RNS_PRIME_BITS'd1110484211, `RNS_PRIME_BITS'd962210911, `RNS_PRIME_BITS'd1051786406, `RNS_PRIME_BITS'd595850019},
    '{`RNS_PRIME_BITS'd1491102736, `RNS_PRIME_BITS'd1997054115, `RNS_PRIME_BITS'd1217383725, `RNS_PRIME_BITS'd744162357, `RNS_PRIME_BITS'd51253230, `RNS_PRIME_BITS'd541786111, `RNS_PRIME_BITS'd1609158059, `RNS_PRIME_BITS'd441302679, `RNS_PRIME_BITS'd1848214536, `RNS_PRIME_BITS'd647462316},
    '{`RNS_PRIME_BITS'd2021134738, `RNS_PRIME_BITS'd794776015, `RNS_PRIME_BITS'd1863885714, `RNS_PRIME_BITS'd1279192758, `RNS_PRIME_BITS'd1485198861, `RNS_PRIME_BITS'd1272035409, `RNS_PRIME_BITS'd720349947, `RNS_PRIME_BITS'd1885474451, `RNS_PRIME_BITS'd531632460, `RNS_PRIME_BITS'd621807479},
    '{`RNS_PRIME_BITS'd1579513695, `RNS_PRIME_BITS'd1314130912, `RNS_PRIME_BITS'd323928954, `RNS_PRIME_BITS'd410212018, `RNS_PRIME_BITS'd233960928, `RNS_PRIME_BITS'd341624221, `RNS_PRIME_BITS'd484991355, `RNS_PRIME_BITS'd1709782841, `RNS_PRIME_BITS'd1716054783, `RNS_PRIME_BITS'd2086146408},
    '{`RNS_PRIME_BITS'd1833484025, `RNS_PRIME_BITS'd973053246, `RNS_PRIME_BITS'd996358001, `RNS_PRIME_BITS'd290057533, `RNS_PRIME_BITS'd1255713559, `RNS_PRIME_BITS'd600566031, `RNS_PRIME_BITS'd97355034, `RNS_PRIME_BITS'd1991992747, `RNS_PRIME_BITS'd1013332612, `RNS_PRIME_BITS'd21134795},
    '{`RNS_PRIME_BITS'd415407688, `RNS_PRIME_BITS'd390565408, `RNS_PRIME_BITS'd1381860284, `RNS_PRIME_BITS'd1950371777, `RNS_PRIME_BITS'd653561290, `RNS_PRIME_BITS'd86629881, `RNS_PRIME_BITS'd1645756096, `RNS_PRIME_BITS'd1105271508, `RNS_PRIME_BITS'd8508976, `RNS_PRIME_BITS'd1095737960},
    '{`RNS_PRIME_BITS'd108410860, `RNS_PRIME_BITS'd2078087010, `RNS_PRIME_BITS'd1957249992, `RNS_PRIME_BITS'd1175837644, `RNS_PRIME_BITS'd1809274866, `RNS_PRIME_BITS'd1340574042, `RNS_PRIME_BITS'd661533370, `RNS_PRIME_BITS'd1959824221, `RNS_PRIME_BITS'd1812041745, `RNS_PRIME_BITS'd1659943279},
    '{`RNS_PRIME_BITS'd390012958, `RNS_PRIME_BITS'd2117437096, `RNS_PRIME_BITS'd409065623, `RNS_PRIME_BITS'd981070349, `RNS_PRIME_BITS'd1291309433, `RNS_PRIME_BITS'd2011139044, `RNS_PRIME_BITS'd732721758, `RNS_PRIME_BITS'd518766479, `RNS_PRIME_BITS'd1294117088, `RNS_PRIME_BITS'd818892796},
    '{`RNS_PRIME_BITS'd39513013, `RNS_PRIME_BITS'd2143795973, `RNS_PRIME_BITS'd1434802343, `RNS_PRIME_BITS'd614980717, `RNS_PRIME_BITS'd1460419000, `RNS_PRIME_BITS'd1086315716, `RNS_PRIME_BITS'd857228700, `RNS_PRIME_BITS'd439717886, `RNS_PRIME_BITS'd602291994, `RNS_PRIME_BITS'd1131234638},
    '{`RNS_PRIME_BITS'd1315307254, `RNS_PRIME_BITS'd690802843, `RNS_PRIME_BITS'd1224672529, `RNS_PRIME_BITS'd579582540, `RNS_PRIME_BITS'd856192602, `RNS_PRIME_BITS'd1531478782, `RNS_PRIME_BITS'd1020718827, `RNS_PRIME_BITS'd709867172, `RNS_PRIME_BITS'd1262688818, `RNS_PRIME_BITS'd737003659},
    '{`RNS_PRIME_BITS'd1035956851, `RNS_PRIME_BITS'd80921750, `RNS_PRIME_BITS'd1715559177, `RNS_PRIME_BITS'd1508357394, `RNS_PRIME_BITS'd1435552928, `RNS_PRIME_BITS'd1539211725, `RNS_PRIME_BITS'd1709935961, `RNS_PRIME_BITS'd699131328, `RNS_PRIME_BITS'd1869509655, `RNS_PRIME_BITS'd152293315},
    '{`RNS_PRIME_BITS'd2147353437, `RNS_PRIME_BITS'd114305354, `RNS_PRIME_BITS'd760603346, `RNS_PRIME_BITS'd1273694749, `RNS_PRIME_BITS'd1935378783, `RNS_PRIME_BITS'd1734988592, `RNS_PRIME_BITS'd431737100, `RNS_PRIME_BITS'd1291524712, `RNS_PRIME_BITS'd1960509946, `RNS_PRIME_BITS'd712173292},
    '{`RNS_PRIME_BITS'd766995009, `RNS_PRIME_BITS'd1165772423, `RNS_PRIME_BITS'd25741449, `RNS_PRIME_BITS'd1914103360, `RNS_PRIME_BITS'd2081438194, `RNS_PRIME_BITS'd1990344641, `RNS_PRIME_BITS'd732679864, `RNS_PRIME_BITS'd774912588, `RNS_PRIME_BITS'd1714061643, `RNS_PRIME_BITS'd840211036},
    '{`RNS_PRIME_BITS'd1736119076, `RNS_PRIME_BITS'd1291865825, `RNS_PRIME_BITS'd1857266219, `RNS_PRIME_BITS'd912129036, `RNS_PRIME_BITS'd1577082940, `RNS_PRIME_BITS'd2057659125, `RNS_PRIME_BITS'd671545775, `RNS_PRIME_BITS'd1483619555, `RNS_PRIME_BITS'd2035490122, `RNS_PRIME_BITS'd701151613},
    '{`RNS_PRIME_BITS'd1671136753, `RNS_PRIME_BITS'd1902067646, `RNS_PRIME_BITS'd802239014, `RNS_PRIME_BITS'd240464665, `RNS_PRIME_BITS'd1248652945, `RNS_PRIME_BITS'd1918694108, `RNS_PRIME_BITS'd1818415756, `RNS_PRIME_BITS'd1717733819, `RNS_PRIME_BITS'd1805451593, `RNS_PRIME_BITS'd1118340653},
    '{`RNS_PRIME_BITS'd1852152637, `RNS_PRIME_BITS'd591989474, `RNS_PRIME_BITS'd1490051286, `RNS_PRIME_BITS'd1828694336, `RNS_PRIME_BITS'd533947106, `RNS_PRIME_BITS'd776836116, `RNS_PRIME_BITS'd266352970, `RNS_PRIME_BITS'd2144615113, `RNS_PRIME_BITS'd480486321, `RNS_PRIME_BITS'd2008388677},
    '{`RNS_PRIME_BITS'd679154017, `RNS_PRIME_BITS'd1358610859, `RNS_PRIME_BITS'd1183045395, `RNS_PRIME_BITS'd1311123035, `RNS_PRIME_BITS'd1859122038, `RNS_PRIME_BITS'd2113226479, `RNS_PRIME_BITS'd34150006, `RNS_PRIME_BITS'd923129522, `RNS_PRIME_BITS'd1348869430, `RNS_PRIME_BITS'd901615418},
    '{`RNS_PRIME_BITS'd1903872203, `RNS_PRIME_BITS'd1213908812, `RNS_PRIME_BITS'd817750688, `RNS_PRIME_BITS'd1470475081, `RNS_PRIME_BITS'd522771328, `RNS_PRIME_BITS'd1619685630, `RNS_PRIME_BITS'd639777332, `RNS_PRIME_BITS'd1782014888, `RNS_PRIME_BITS'd210379497, `RNS_PRIME_BITS'd1631682801},
    '{`RNS_PRIME_BITS'd509803209, `RNS_PRIME_BITS'd1456157157, `RNS_PRIME_BITS'd452894477, `RNS_PRIME_BITS'd1947779633, `RNS_PRIME_BITS'd406008748, `RNS_PRIME_BITS'd1532292834, `RNS_PRIME_BITS'd1994110563, `RNS_PRIME_BITS'd498329367, `RNS_PRIME_BITS'd219162379, `RNS_PRIME_BITS'd894989546},
    '{`RNS_PRIME_BITS'd1923228553, `RNS_PRIME_BITS'd1512379339, `RNS_PRIME_BITS'd1795586742, `RNS_PRIME_BITS'd1907459693, `RNS_PRIME_BITS'd438860140, `RNS_PRIME_BITS'd1701484285, `RNS_PRIME_BITS'd17290594, `RNS_PRIME_BITS'd1916044635, `RNS_PRIME_BITS'd1148913620, `RNS_PRIME_BITS'd1219619620},
    '{`RNS_PRIME_BITS'd2117832527, `RNS_PRIME_BITS'd815983636, `RNS_PRIME_BITS'd961636590, `RNS_PRIME_BITS'd658894168, `RNS_PRIME_BITS'd1210778163, `RNS_PRIME_BITS'd2119146802, `RNS_PRIME_BITS'd701266969, `RNS_PRIME_BITS'd1266466375, `RNS_PRIME_BITS'd305150941, `RNS_PRIME_BITS'd181570311},
    '{`RNS_PRIME_BITS'd1506837361, `RNS_PRIME_BITS'd88552478, `RNS_PRIME_BITS'd933771280, `RNS_PRIME_BITS'd241969214, `RNS_PRIME_BITS'd489034685, `RNS_PRIME_BITS'd1774678146, `RNS_PRIME_BITS'd389917424, `RNS_PRIME_BITS'd1566242377, `RNS_PRIME_BITS'd1397283234, `RNS_PRIME_BITS'd865222540},
    '{`RNS_PRIME_BITS'd2079579615, `RNS_PRIME_BITS'd1971063340, `RNS_PRIME_BITS'd2067250763, `RNS_PRIME_BITS'd1268920098, `RNS_PRIME_BITS'd418699502, `RNS_PRIME_BITS'd1965954990, `RNS_PRIME_BITS'd526726797, `RNS_PRIME_BITS'd413468582, `RNS_PRIME_BITS'd2006122730, `RNS_PRIME_BITS'd1450038462},
    '{`RNS_PRIME_BITS'd1250823470, `RNS_PRIME_BITS'd1752621452, `RNS_PRIME_BITS'd1606867391, `RNS_PRIME_BITS'd1482500299, `RNS_PRIME_BITS'd762464778, `RNS_PRIME_BITS'd252985111, `RNS_PRIME_BITS'd2045270253, `RNS_PRIME_BITS'd643788293, `RNS_PRIME_BITS'd171919279, `RNS_PRIME_BITS'd1234398263},
    '{`RNS_PRIME_BITS'd420228658, `RNS_PRIME_BITS'd1862643389, `RNS_PRIME_BITS'd1587391278, `RNS_PRIME_BITS'd2139683486, `RNS_PRIME_BITS'd2015785457, `RNS_PRIME_BITS'd1613231448, `RNS_PRIME_BITS'd494146855, `RNS_PRIME_BITS'd1094515363, `RNS_PRIME_BITS'd536327602, `RNS_PRIME_BITS'd823293093},
    '{`RNS_PRIME_BITS'd1563075904, `RNS_PRIME_BITS'd1172681457, `RNS_PRIME_BITS'd1867891810, `RNS_PRIME_BITS'd182401501, `RNS_PRIME_BITS'd82736443, `RNS_PRIME_BITS'd1791618311, `RNS_PRIME_BITS'd51676344, `RNS_PRIME_BITS'd1240667604, `RNS_PRIME_BITS'd1329388365, `RNS_PRIME_BITS'd1985363596},
    '{`RNS_PRIME_BITS'd502881983, `RNS_PRIME_BITS'd1143682806, `RNS_PRIME_BITS'd791946393, `RNS_PRIME_BITS'd404297573, `RNS_PRIME_BITS'd1147732095, `RNS_PRIME_BITS'd1019893963, `RNS_PRIME_BITS'd1682210285, `RNS_PRIME_BITS'd543457931, `RNS_PRIME_BITS'd1974613206, `RNS_PRIME_BITS'd818331108},
    '{`RNS_PRIME_BITS'd724031645, `RNS_PRIME_BITS'd338550976, `RNS_PRIME_BITS'd1977528817, `RNS_PRIME_BITS'd600086169, `RNS_PRIME_BITS'd1784510466, `RNS_PRIME_BITS'd656790317, `RNS_PRIME_BITS'd11799338, `RNS_PRIME_BITS'd1937502361, `RNS_PRIME_BITS'd676472523, `RNS_PRIME_BITS'd1561855482},
    '{`RNS_PRIME_BITS'd1772628239, `RNS_PRIME_BITS'd106453541, `RNS_PRIME_BITS'd1333056578, `RNS_PRIME_BITS'd1898969837, `RNS_PRIME_BITS'd616269263, `RNS_PRIME_BITS'd2095773699, `RNS_PRIME_BITS'd605994818, `RNS_PRIME_BITS'd302758082, `RNS_PRIME_BITS'd516841753, `RNS_PRIME_BITS'd1162473475},
    '{`RNS_PRIME_BITS'd1192992316, `RNS_PRIME_BITS'd2025614866, `RNS_PRIME_BITS'd1936618199, `RNS_PRIME_BITS'd381798226, `RNS_PRIME_BITS'd1568211351, `RNS_PRIME_BITS'd475509346, `RNS_PRIME_BITS'd810520533, `RNS_PRIME_BITS'd1245689600, `RNS_PRIME_BITS'd1635059530, `RNS_PRIME_BITS'd679665385},
    '{`RNS_PRIME_BITS'd799510527, `RNS_PRIME_BITS'd1520721165, `RNS_PRIME_BITS'd394575869, `RNS_PRIME_BITS'd1471656364, `RNS_PRIME_BITS'd996647107, `RNS_PRIME_BITS'd1766991867, `RNS_PRIME_BITS'd466318405, `RNS_PRIME_BITS'd233735314, `RNS_PRIME_BITS'd206088228, `RNS_PRIME_BITS'd151684780},
    '{`RNS_PRIME_BITS'd865281393, `RNS_PRIME_BITS'd451495488, `RNS_PRIME_BITS'd1706183883, `RNS_PRIME_BITS'd1883030321, `RNS_PRIME_BITS'd93069258, `RNS_PRIME_BITS'd744474398, `RNS_PRIME_BITS'd1696380915, `RNS_PRIME_BITS'd1244502731, `RNS_PRIME_BITS'd1978964303, `RNS_PRIME_BITS'd189652214},
    '{`RNS_PRIME_BITS'd1440919025, `RNS_PRIME_BITS'd1439260276, `RNS_PRIME_BITS'd1019994178, `RNS_PRIME_BITS'd1910553218, `RNS_PRIME_BITS'd109889889, `RNS_PRIME_BITS'd1385528499, `RNS_PRIME_BITS'd1411989176, `RNS_PRIME_BITS'd417947728, `RNS_PRIME_BITS'd530277962, `RNS_PRIME_BITS'd368403599},
    '{`RNS_PRIME_BITS'd320919212, `RNS_PRIME_BITS'd470089507, `RNS_PRIME_BITS'd2110959079, `RNS_PRIME_BITS'd560223679, `RNS_PRIME_BITS'd1857149402, `RNS_PRIME_BITS'd1683141286, `RNS_PRIME_BITS'd691036032, `RNS_PRIME_BITS'd1315190558, `RNS_PRIME_BITS'd518870814, `RNS_PRIME_BITS'd1529671476},
    '{`RNS_PRIME_BITS'd1425746572, `RNS_PRIME_BITS'd1915228943, `RNS_PRIME_BITS'd448377474, `RNS_PRIME_BITS'd1314210880, `RNS_PRIME_BITS'd134831017, `RNS_PRIME_BITS'd789157594, `RNS_PRIME_BITS'd262413762, `RNS_PRIME_BITS'd387463468, `RNS_PRIME_BITS'd1100050078, `RNS_PRIME_BITS'd1835710782},
    '{`RNS_PRIME_BITS'd194388085, `RNS_PRIME_BITS'd1497132433, `RNS_PRIME_BITS'd405699713, `RNS_PRIME_BITS'd773746588, `RNS_PRIME_BITS'd1147529730, `RNS_PRIME_BITS'd709285475, `RNS_PRIME_BITS'd796850585, `RNS_PRIME_BITS'd8513528, `RNS_PRIME_BITS'd1223389601, `RNS_PRIME_BITS'd809821929},
    '{`RNS_PRIME_BITS'd1911050575, `RNS_PRIME_BITS'd1272580642, `RNS_PRIME_BITS'd1086763977, `RNS_PRIME_BITS'd1879403728, `RNS_PRIME_BITS'd1866444078, `RNS_PRIME_BITS'd1679060775, `RNS_PRIME_BITS'd213096340, `RNS_PRIME_BITS'd363824824, `RNS_PRIME_BITS'd232806416, `RNS_PRIME_BITS'd1467187245},
    '{`RNS_PRIME_BITS'd157744050, `RNS_PRIME_BITS'd317748997, `RNS_PRIME_BITS'd949740882, `RNS_PRIME_BITS'd857339974, `RNS_PRIME_BITS'd2144032563, `RNS_PRIME_BITS'd1793260831, `RNS_PRIME_BITS'd1262742624, `RNS_PRIME_BITS'd714600989, `RNS_PRIME_BITS'd2109715245, `RNS_PRIME_BITS'd534996762},
    '{`RNS_PRIME_BITS'd364446835, `RNS_PRIME_BITS'd640153685, `RNS_PRIME_BITS'd1548919159, `RNS_PRIME_BITS'd137873604, `RNS_PRIME_BITS'd55494586, `RNS_PRIME_BITS'd219448318, `RNS_PRIME_BITS'd1034174435, `RNS_PRIME_BITS'd908083776, `RNS_PRIME_BITS'd1009260182, `RNS_PRIME_BITS'd562322150},
    '{`RNS_PRIME_BITS'd814191722, `RNS_PRIME_BITS'd2014711680, `RNS_PRIME_BITS'd2103401360, `RNS_PRIME_BITS'd945427192, `RNS_PRIME_BITS'd680948919, `RNS_PRIME_BITS'd1848718917, `RNS_PRIME_BITS'd854251826, `RNS_PRIME_BITS'd352065477, `RNS_PRIME_BITS'd1880309153, `RNS_PRIME_BITS'd2032895388},
    '{`RNS_PRIME_BITS'd294646135, `RNS_PRIME_BITS'd858062951, `RNS_PRIME_BITS'd382100498, `RNS_PRIME_BITS'd1095830114, `RNS_PRIME_BITS'd327764410, `RNS_PRIME_BITS'd192946793, `RNS_PRIME_BITS'd1299115799, `RNS_PRIME_BITS'd135517024, `RNS_PRIME_BITS'd255993234, `RNS_PRIME_BITS'd791949256},
    '{`RNS_PRIME_BITS'd1813437066, `RNS_PRIME_BITS'd1376521486, `RNS_PRIME_BITS'd921953420, `RNS_PRIME_BITS'd1623445789, `RNS_PRIME_BITS'd1002175446, `RNS_PRIME_BITS'd637515552, `RNS_PRIME_BITS'd1227114396, `RNS_PRIME_BITS'd929671741, `RNS_PRIME_BITS'd73643954, `RNS_PRIME_BITS'd1077481907},
    '{`RNS_PRIME_BITS'd1157933193, `RNS_PRIME_BITS'd588621655, `RNS_PRIME_BITS'd2104639994, `RNS_PRIME_BITS'd754910642, `RNS_PRIME_BITS'd679940496, `RNS_PRIME_BITS'd1472261172, `RNS_PRIME_BITS'd1205424420, `RNS_PRIME_BITS'd1955644931, `RNS_PRIME_BITS'd365178688, `RNS_PRIME_BITS'd1194674271},
    '{`RNS_PRIME_BITS'd581524369, `RNS_PRIME_BITS'd1400761654, `RNS_PRIME_BITS'd453375438, `RNS_PRIME_BITS'd372240821, `RNS_PRIME_BITS'd1943465816, `RNS_PRIME_BITS'd2129800416, `RNS_PRIME_BITS'd1374254703, `RNS_PRIME_BITS'd1084106769, `RNS_PRIME_BITS'd1687722945, `RNS_PRIME_BITS'd381452777},
    '{`RNS_PRIME_BITS'd1043594109, `RNS_PRIME_BITS'd1475140116, `RNS_PRIME_BITS'd989282524, `RNS_PRIME_BITS'd1883104327, `RNS_PRIME_BITS'd1565393479, `RNS_PRIME_BITS'd1358992016, `RNS_PRIME_BITS'd2061921710, `RNS_PRIME_BITS'd1211141776, `RNS_PRIME_BITS'd1194694038, `RNS_PRIME_BITS'd2104040240},
    '{`RNS_PRIME_BITS'd2040809068, `RNS_PRIME_BITS'd2044949706, `RNS_PRIME_BITS'd1935554307, `RNS_PRIME_BITS'd1666316763, `RNS_PRIME_BITS'd723203597, `RNS_PRIME_BITS'd281731676, `RNS_PRIME_BITS'd925175951, `RNS_PRIME_BITS'd431309378, `RNS_PRIME_BITS'd1089849203, `RNS_PRIME_BITS'd197504372},
    '{`RNS_PRIME_BITS'd1362467077, `RNS_PRIME_BITS'd369013195, `RNS_PRIME_BITS'd147736310, `RNS_PRIME_BITS'd436763432, `RNS_PRIME_BITS'd296932084, `RNS_PRIME_BITS'd351224846, `RNS_PRIME_BITS'd1059549025, `RNS_PRIME_BITS'd1448015126, `RNS_PRIME_BITS'd710114276, `RNS_PRIME_BITS'd945201478},
    '{`RNS_PRIME_BITS'd1840385618, `RNS_PRIME_BITS'd239274132, `RNS_PRIME_BITS'd1380723173, `RNS_PRIME_BITS'd980861161, `RNS_PRIME_BITS'd1471067818, `RNS_PRIME_BITS'd1440309923, `RNS_PRIME_BITS'd130866692, `RNS_PRIME_BITS'd580446224, `RNS_PRIME_BITS'd586395470, `RNS_PRIME_BITS'd1372404310},
    '{`RNS_PRIME_BITS'd786034799, `RNS_PRIME_BITS'd1369478611, `RNS_PRIME_BITS'd426314629, `RNS_PRIME_BITS'd898924278, `RNS_PRIME_BITS'd483249824, `RNS_PRIME_BITS'd1372906079, `RNS_PRIME_BITS'd212330703, `RNS_PRIME_BITS'd598644579, `RNS_PRIME_BITS'd533019697, `RNS_PRIME_BITS'd1194991604},
    '{`RNS_PRIME_BITS'd1290751872, `RNS_PRIME_BITS'd2121640298, `RNS_PRIME_BITS'd675455857, `RNS_PRIME_BITS'd739943696, `RNS_PRIME_BITS'd2118967517, `RNS_PRIME_BITS'd724776185, `RNS_PRIME_BITS'd1961743338, `RNS_PRIME_BITS'd1344324524, `RNS_PRIME_BITS'd785507157, `RNS_PRIME_BITS'd1695765452},
    '{`RNS_PRIME_BITS'd1835299179, `RNS_PRIME_BITS'd178973199, `RNS_PRIME_BITS'd192169418, `RNS_PRIME_BITS'd1179634056, `RNS_PRIME_BITS'd1906177344, `RNS_PRIME_BITS'd2007997618, `RNS_PRIME_BITS'd1420586335, `RNS_PRIME_BITS'd1710872373, `RNS_PRIME_BITS'd944229547, `RNS_PRIME_BITS'd1967628692},
    '{`RNS_PRIME_BITS'd921535806, `RNS_PRIME_BITS'd1530938706, `RNS_PRIME_BITS'd2075195857, `RNS_PRIME_BITS'd1871358114, `RNS_PRIME_BITS'd1709697570, `RNS_PRIME_BITS'd373483603, `RNS_PRIME_BITS'd1451380014, `RNS_PRIME_BITS'd2029814002, `RNS_PRIME_BITS'd621626299, `RNS_PRIME_BITS'd113472302},
    '{`RNS_PRIME_BITS'd1736524985, `RNS_PRIME_BITS'd851381315, `RNS_PRIME_BITS'd794958276, `RNS_PRIME_BITS'd1686287107, `RNS_PRIME_BITS'd471423405, `RNS_PRIME_BITS'd1314350158, `RNS_PRIME_BITS'd1356634446, `RNS_PRIME_BITS'd997666869, `RNS_PRIME_BITS'd282182630, `RNS_PRIME_BITS'd367143186},
    '{`RNS_PRIME_BITS'd1772903848, `RNS_PRIME_BITS'd473394055, `RNS_PRIME_BITS'd517015927, `RNS_PRIME_BITS'd1063638444, `RNS_PRIME_BITS'd1151883039, `RNS_PRIME_BITS'd1924854916, `RNS_PRIME_BITS'd1147962701, `RNS_PRIME_BITS'd1393964494, `RNS_PRIME_BITS'd1181715581, `RNS_PRIME_BITS'd113949623},
    '{`RNS_PRIME_BITS'd1639441736, `RNS_PRIME_BITS'd1892140015, `RNS_PRIME_BITS'd472050077, `RNS_PRIME_BITS'd257841232, `RNS_PRIME_BITS'd1176332907, `RNS_PRIME_BITS'd231705128, `RNS_PRIME_BITS'd1856735785, `RNS_PRIME_BITS'd1467479091, `RNS_PRIME_BITS'd233193577, `RNS_PRIME_BITS'd1307104724},
    '{`RNS_PRIME_BITS'd875963076, `RNS_PRIME_BITS'd545148602, `RNS_PRIME_BITS'd793838922, `RNS_PRIME_BITS'd1619378277, `RNS_PRIME_BITS'd1142358308, `RNS_PRIME_BITS'd882304718, `RNS_PRIME_BITS'd1296291999, `RNS_PRIME_BITS'd93058891, `RNS_PRIME_BITS'd1167177632, `RNS_PRIME_BITS'd1811708202},
    '{`RNS_PRIME_BITS'd631964093, `RNS_PRIME_BITS'd1078734864, `RNS_PRIME_BITS'd1410940662, `RNS_PRIME_BITS'd931215593, `RNS_PRIME_BITS'd143724095, `RNS_PRIME_BITS'd1715120914, `RNS_PRIME_BITS'd145347728, `RNS_PRIME_BITS'd377262823, `RNS_PRIME_BITS'd327707007, `RNS_PRIME_BITS'd936229520},
    '{`RNS_PRIME_BITS'd1737368185, `RNS_PRIME_BITS'd111736972, `RNS_PRIME_BITS'd775107127, `RNS_PRIME_BITS'd128280690, `RNS_PRIME_BITS'd1806198909, `RNS_PRIME_BITS'd1907790616, `RNS_PRIME_BITS'd46582280, `RNS_PRIME_BITS'd796221513, `RNS_PRIME_BITS'd1982229971, `RNS_PRIME_BITS'd118485329},
    '{`RNS_PRIME_BITS'd443906989, `RNS_PRIME_BITS'd1874084926, `RNS_PRIME_BITS'd1905445759, `RNS_PRIME_BITS'd1249145541, `RNS_PRIME_BITS'd1372271781, `RNS_PRIME_BITS'd709800044, `RNS_PRIME_BITS'd1151694911, `RNS_PRIME_BITS'd587837481, `RNS_PRIME_BITS'd614945244, `RNS_PRIME_BITS'd733045511},
    '{`RNS_PRIME_BITS'd420854524, `RNS_PRIME_BITS'd1635406236, `RNS_PRIME_BITS'd1827960, `RNS_PRIME_BITS'd595856712, `RNS_PRIME_BITS'd641242964, `RNS_PRIME_BITS'd1861693614, `RNS_PRIME_BITS'd2126926337, `RNS_PRIME_BITS'd268706943, `RNS_PRIME_BITS'd1143589008, `RNS_PRIME_BITS'd91268120}
};

parameter Ba_BASIS_poly twist_factor_ba   = '{
    '{`RNS_PRIME_BITS'd1},
    '{`RNS_PRIME_BITS'd408088301},
    '{`RNS_PRIME_BITS'd545722081},
    '{`RNS_PRIME_BITS'd2013316613},
    '{`RNS_PRIME_BITS'd1321642193},
    '{`RNS_PRIME_BITS'd321959319},
    '{`RNS_PRIME_BITS'd1021511790},
    '{`RNS_PRIME_BITS'd895733675},
    '{`RNS_PRIME_BITS'd1907272939},
    '{`RNS_PRIME_BITS'd1047887518},
    '{`RNS_PRIME_BITS'd130472541},
    '{`RNS_PRIME_BITS'd849014309},
    '{`RNS_PRIME_BITS'd1383024311},
    '{`RNS_PRIME_BITS'd2051297149},
    '{`RNS_PRIME_BITS'd572408039},
    '{`RNS_PRIME_BITS'd708487692},
    '{`RNS_PRIME_BITS'd1187016878},
    '{`RNS_PRIME_BITS'd1217688897},
    '{`RNS_PRIME_BITS'd1748729974},
    '{`RNS_PRIME_BITS'd1671387385},
    '{`RNS_PRIME_BITS'd2040483268},
    '{`RNS_PRIME_BITS'd985132875},
    '{`RNS_PRIME_BITS'd1013309155},
    '{`RNS_PRIME_BITS'd1103304400},
    '{`RNS_PRIME_BITS'd70525087},
    '{`RNS_PRIME_BITS'd1280246740},
    '{`RNS_PRIME_BITS'd1423738182},
    '{`RNS_PRIME_BITS'd2108544873},
    '{`RNS_PRIME_BITS'd1332271570},
    '{`RNS_PRIME_BITS'd1752678097},
    '{`RNS_PRIME_BITS'd658442757},
    '{`RNS_PRIME_BITS'd427090976},
    '{`RNS_PRIME_BITS'd1656931938},
    '{`RNS_PRIME_BITS'd828187205},
    '{`RNS_PRIME_BITS'd863028180},
    '{`RNS_PRIME_BITS'd1908486966},
    '{`RNS_PRIME_BITS'd61269856},
    '{`RNS_PRIME_BITS'd1612421805},
    '{`RNS_PRIME_BITS'd1825676708},
    '{`RNS_PRIME_BITS'd1310355683},
    '{`RNS_PRIME_BITS'd99928383},
    '{`RNS_PRIME_BITS'd1003955160},
    '{`RNS_PRIME_BITS'd1348001053},
    '{`RNS_PRIME_BITS'd819422651},
    '{`RNS_PRIME_BITS'd1070648195},
    '{`RNS_PRIME_BITS'd1226417430},
    '{`RNS_PRIME_BITS'd1453801843},
    '{`RNS_PRIME_BITS'd997812037},
    '{`RNS_PRIME_BITS'd163057938},
    '{`RNS_PRIME_BITS'd583652742},
    '{`RNS_PRIME_BITS'd1898138826},
    '{`RNS_PRIME_BITS'd1278600277},
    '{`RNS_PRIME_BITS'd1437033183},
    '{`RNS_PRIME_BITS'd2058685992},
    '{`RNS_PRIME_BITS'd2047246327},
    '{`RNS_PRIME_BITS'd2003019592},
    '{`RNS_PRIME_BITS'd608435798},
    '{`RNS_PRIME_BITS'd843307226},
    '{`RNS_PRIME_BITS'd881750696},
    '{`RNS_PRIME_BITS'd52620857},
    '{`RNS_PRIME_BITS'd1434548924},
    '{`RNS_PRIME_BITS'd618722642},
    '{`RNS_PRIME_BITS'd1713622070},
    '{`RNS_PRIME_BITS'd2138310495}
};

parameter Ba_BASIS_poly untwist_factor_ba = '{
    '{`RNS_PRIME_BITS'd2113948747},
    '{`RNS_PRIME_BITS'd1006785901},
    '{`RNS_PRIME_BITS'd1785180724},
    '{`RNS_PRIME_BITS'd594317815},
    '{`RNS_PRIME_BITS'd1990869694},
    '{`RNS_PRIME_BITS'd1911798094},
    '{`RNS_PRIME_BITS'd1328412326},
    '{`RNS_PRIME_BITS'd859246617},
    '{`RNS_PRIME_BITS'd728697515},
    '{`RNS_PRIME_BITS'd237140755},
    '{`RNS_PRIME_BITS'd1813522587},
    '{`RNS_PRIME_BITS'd1310022712},
    '{`RNS_PRIME_BITS'd1017743359},
    '{`RNS_PRIME_BITS'd684671453},
    '{`RNS_PRIME_BITS'd305889001},
    '{`RNS_PRIME_BITS'd192208878},
    '{`RNS_PRIME_BITS'd601437576},
    '{`RNS_PRIME_BITS'd152182897},
    '{`RNS_PRIME_BITS'd1688576189},
    '{`RNS_PRIME_BITS'd719041552},
    '{`RNS_PRIME_BITS'd83935348},
    '{`RNS_PRIME_BITS'd1966926300},
    '{`RNS_PRIME_BITS'd952025002},
    '{`RNS_PRIME_BITS'd789627009},
    '{`RNS_PRIME_BITS'd2112387366},
    '{`RNS_PRIME_BITS'd1153941663},
    '{`RNS_PRIME_BITS'd1179444514},
    '{`RNS_PRIME_BITS'd1484769300},
    '{`RNS_PRIME_BITS'd1072794403},
    '{`RNS_PRIME_BITS'd1782135960},
    '{`RNS_PRIME_BITS'd657610025},
    '{`RNS_PRIME_BITS'd154833285},
    '{`RNS_PRIME_BITS'd1114971667},
    '{`RNS_PRIME_BITS'd1067078448},
    '{`RNS_PRIME_BITS'd157485542},
    '{`RNS_PRIME_BITS'd543045019},
    '{`RNS_PRIME_BITS'd583168613},
    '{`RNS_PRIME_BITS'd1342798409},
    '{`RNS_PRIME_BITS'd179082543},
    '{`RNS_PRIME_BITS'd651090985},
    '{`RNS_PRIME_BITS'd1039095048},
    '{`RNS_PRIME_BITS'd519636741},
    '{`RNS_PRIME_BITS'd1158583015},
    '{`RNS_PRIME_BITS'd353709461},
    '{`RNS_PRIME_BITS'd102336417},
    '{`RNS_PRIME_BITS'd1886504867},
    '{`RNS_PRIME_BITS'd1784632163},
    '{`RNS_PRIME_BITS'd14528353},
    '{`RNS_PRIME_BITS'd1524970994},
    '{`RNS_PRIME_BITS'd391586784},
    '{`RNS_PRIME_BITS'd1299691063},
    '{`RNS_PRIME_BITS'd2014787745},
    '{`RNS_PRIME_BITS'd1823901056},
    '{`RNS_PRIME_BITS'd1228259606},
    '{`RNS_PRIME_BITS'd971048885},
    '{`RNS_PRIME_BITS'd990269018},
    '{`RNS_PRIME_BITS'd1413052767},
    '{`RNS_PRIME_BITS'd1428858068},
    '{`RNS_PRIME_BITS'd1527557011},
    '{`RNS_PRIME_BITS'd766728452},
    '{`RNS_PRIME_BITS'd549779955},
    '{`RNS_PRIME_BITS'd136315638},
    '{`RNS_PRIME_BITS'd1098779579},
    '{`RNS_PRIME_BITS'd1503587011}
};


// fastBConv precalculated inverses
parameter rns_residue_t z_MOD_q[`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1340848717, `RNS_PRIME_BITS'd1950706637, `RNS_PRIME_BITS'd136505383, `RNS_PRIME_BITS'd1261863396, `RNS_PRIME_BITS'd490720514, `RNS_PRIME_BITS'd2048232271, `RNS_PRIME_BITS'd561180295, `RNS_PRIME_BITS'd2064343317, `RNS_PRIME_BITS'd1284162414, `RNS_PRIME_BITS'd426116969};
parameter rns_residue_t z_MOD_B[`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd400603566, `RNS_PRIME_BITS'd1317047788, `RNS_PRIME_BITS'd1877527982, `RNS_PRIME_BITS'd816591707, `RNS_PRIME_BITS'd1500256234, `RNS_PRIME_BITS'd8640588, `RNS_PRIME_BITS'd1509953789, `RNS_PRIME_BITS'd1256593971, `RNS_PRIME_BITS'd1660146682, `RNS_PRIME_BITS'd390117507};
parameter rns_residue_t y_q_TO_qBBa[`qBBa_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1514938357, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1663002026, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1202970911, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1254269319, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd15070697, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd93592423, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd345241794, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd126359634, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1571891470, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1004678308 },
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};
parameter rns_residue_t y_B_TO_Ba[`Ba_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd33728781, `RNS_PRIME_BITS'd1756228743, `RNS_PRIME_BITS'd487215260, `RNS_PRIME_BITS'd501135696, `RNS_PRIME_BITS'd459470026, `RNS_PRIME_BITS'd1877657833, `RNS_PRIME_BITS'd50297305, `RNS_PRIME_BITS'd56214635, `RNS_PRIME_BITS'd1200871039, `RNS_PRIME_BITS'd1750218591 }
};
parameter rns_residue_t y_B_TO_q[`q_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd10, `RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd92 },
'{ `RNS_PRIME_BITS'd1219156511, `RNS_PRIME_BITS'd1608499681, `RNS_PRIME_BITS'd371154937, `RNS_PRIME_BITS'd924754142, `RNS_PRIME_BITS'd2003633539, `RNS_PRIME_BITS'd627440795, `RNS_PRIME_BITS'd1066486116, `RNS_PRIME_BITS'd1296251710, `RNS_PRIME_BITS'd1679092476, `RNS_PRIME_BITS'd772683368 },
'{ `RNS_PRIME_BITS'd1367502590, `RNS_PRIME_BITS'd1413619003, `RNS_PRIME_BITS'd1604587363, `RNS_PRIME_BITS'd796115568, `RNS_PRIME_BITS'd154115966, `RNS_PRIME_BITS'd287007179, `RNS_PRIME_BITS'd457558717, `RNS_PRIME_BITS'd43558045, `RNS_PRIME_BITS'd1825868505, `RNS_PRIME_BITS'd2117666329 },
'{ `RNS_PRIME_BITS'd488607457, `RNS_PRIME_BITS'd725589953, `RNS_PRIME_BITS'd166254356, `RNS_PRIME_BITS'd1679376923, `RNS_PRIME_BITS'd375851890, `RNS_PRIME_BITS'd962572449, `RNS_PRIME_BITS'd40302594, `RNS_PRIME_BITS'd37730088, `RNS_PRIME_BITS'd1726493613, `RNS_PRIME_BITS'd1162981935 },
'{ `RNS_PRIME_BITS'd317361695, `RNS_PRIME_BITS'd1920884754, `RNS_PRIME_BITS'd1303976625, `RNS_PRIME_BITS'd107931280, `RNS_PRIME_BITS'd1804980561, `RNS_PRIME_BITS'd1467513527, `RNS_PRIME_BITS'd1597511531, `RNS_PRIME_BITS'd1771541117, `RNS_PRIME_BITS'd2104139963, `RNS_PRIME_BITS'd695454200 },
'{ `RNS_PRIME_BITS'd875545508, `RNS_PRIME_BITS'd1106807570, `RNS_PRIME_BITS'd531200008, `RNS_PRIME_BITS'd656659131, `RNS_PRIME_BITS'd318605813, `RNS_PRIME_BITS'd571007940, `RNS_PRIME_BITS'd1098654767, `RNS_PRIME_BITS'd1477330056, `RNS_PRIME_BITS'd1569331694, `RNS_PRIME_BITS'd503094350 },
'{ `RNS_PRIME_BITS'd2014745094, `RNS_PRIME_BITS'd1203280856, `RNS_PRIME_BITS'd1874657457, `RNS_PRIME_BITS'd664236066, `RNS_PRIME_BITS'd1343163396, `RNS_PRIME_BITS'd349851856, `RNS_PRIME_BITS'd327986115, `RNS_PRIME_BITS'd1527009020, `RNS_PRIME_BITS'd1664893238, `RNS_PRIME_BITS'd2028124638 },
'{ `RNS_PRIME_BITS'd17214643, `RNS_PRIME_BITS'd1528026480, `RNS_PRIME_BITS'd707649348, `RNS_PRIME_BITS'd506168135, `RNS_PRIME_BITS'd623405378, `RNS_PRIME_BITS'd1082352090, `RNS_PRIME_BITS'd1990243254, `RNS_PRIME_BITS'd747636934, `RNS_PRIME_BITS'd1326828836, `RNS_PRIME_BITS'd1378524818 },
'{ `RNS_PRIME_BITS'd1873007184, `RNS_PRIME_BITS'd1982800586, `RNS_PRIME_BITS'd1616965474, `RNS_PRIME_BITS'd936503592, `RNS_PRIME_BITS'd265687623, `RNS_PRIME_BITS'd555195787, `RNS_PRIME_BITS'd703316243, `RNS_PRIME_BITS'd1230764655, `RNS_PRIME_BITS'd220437154, `RNS_PRIME_BITS'd1158294204 },
'{ `RNS_PRIME_BITS'd1171115647, `RNS_PRIME_BITS'd1636056387, `RNS_PRIME_BITS'd89367338, `RNS_PRIME_BITS'd1569217605, `RNS_PRIME_BITS'd148010597, `RNS_PRIME_BITS'd552135592, `RNS_PRIME_BITS'd1046145070, `RNS_PRIME_BITS'd1622489461, `RNS_PRIME_BITS'd627687042, `RNS_PRIME_BITS'd765167266 },
'{ `RNS_PRIME_BITS'd1810327907, `RNS_PRIME_BITS'd659636710, `RNS_PRIME_BITS'd527709368, `RNS_PRIME_BITS'd1981502868, `RNS_PRIME_BITS'd395782026, `RNS_PRIME_BITS'd1625981468, `RNS_PRIME_BITS'd263854684, `RNS_PRIME_BITS'd1651540472, `RNS_PRIME_BITS'd1368489211, `RNS_PRIME_BITS'd1257824607 }
};
parameter rns_residue_t y_q_TO_BBa[`B_BASIS_LEN +`Ba_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};

// mod switch from qBBa to BBa (precalculated finv constants)
parameter rns_residue_t qinv_MOD_BBa[`BBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd1685594561, `RNS_PRIME_BITS'd1127635584, `RNS_PRIME_BITS'd1831397647, `RNS_PRIME_BITS'd1452117633, `RNS_PRIME_BITS'd1199363927, `RNS_PRIME_BITS'd1821452128, `RNS_PRIME_BITS'd953961963, `RNS_PRIME_BITS'd7988901, `RNS_PRIME_BITS'd645938236, `RNS_PRIME_BITS'd541478048, `RNS_PRIME_BITS'd433791376};

// FastBConvEx precalculated values
parameter logic signed [`RNS_PRIME_BITS-1:0] signed_intb_MOD_q[`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd106647274, `RNS_PRIME_BITS'd1344578301, `RNS_PRIME_BITS'd849098797, `RNS_PRIME_BITS'd122197028, `RNS_PRIME_BITS'd843004628, `RNS_PRIME_BITS'd354764829, `RNS_PRIME_BITS'd1343634408, `RNS_PRIME_BITS'd1274379894, `RNS_PRIME_BITS'd1805079809, `RNS_PRIME_BITS'd1733088297};
parameter rns_residue_t binv_Ba_MOD_Ba[`Ba_BASIS_LEN] = '{ `RNS_PRIME_BITS'd223873475 };


// RLev keys consist of 22 polynomials: 11 primes in the q basis * 2 Rlev keys per prime (one for A one for B)
parameter q_BASIS_poly RL_EVAL_KEYS[`q_BASIS_LEN][2] = '{
	'{
		'{
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd1016656020, `RNS_PRIME_BITS'd1117264220, `RNS_PRIME_BITS'd1959205716, `RNS_PRIME_BITS'd1664904101, `RNS_PRIME_BITS'd1027986276, `RNS_PRIME_BITS'd249673108, `RNS_PRIME_BITS'd899404479, `RNS_PRIME_BITS'd993657939, `RNS_PRIME_BITS'd1645355725, `RNS_PRIME_BITS'd643096553},
			'{`RNS_PRIME_BITS'd40, `RNS_PRIME_BITS'd1156180647, `RNS_PRIME_BITS'd624971294, `RNS_PRIME_BITS'd2092241288, `RNS_PRIME_BITS'd107813485, `RNS_PRIME_BITS'd1918690432, `RNS_PRIME_BITS'd427151719, `RNS_PRIME_BITS'd1110879368, `RNS_PRIME_BITS'd797105280, `RNS_PRIME_BITS'd317357199, `RNS_PRIME_BITS'd1148174967},
			'{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd653150916, `RNS_PRIME_BITS'd1162281652, `RNS_PRIME_BITS'd1900554648, `RNS_PRIME_BITS'd1803990456, `RNS_PRIME_BITS'd746968738, `RNS_PRIME_BITS'd1551584092, `RNS_PRIME_BITS'd2113458810, `RNS_PRIME_BITS'd1742119537, `RNS_PRIME_BITS'd1968061038, `RNS_PRIME_BITS'd2008153718},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd1524174465, `RNS_PRIME_BITS'd1633824692, `RNS_PRIME_BITS'd239018344, `RNS_PRIME_BITS'd457532961, `RNS_PRIME_BITS'd47853266, `RNS_PRIME_BITS'd1134897370, `RNS_PRIME_BITS'd2115139363, `RNS_PRIME_BITS'd1510015780, `RNS_PRIME_BITS'd2036065412, `RNS_PRIME_BITS'd2049241068},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1402855555, `RNS_PRIME_BITS'd476428980, `RNS_PRIME_BITS'd493392748, `RNS_PRIME_BITS'd1069479952, `RNS_PRIME_BITS'd36577808, `RNS_PRIME_BITS'd247912784, `RNS_PRIME_BITS'd326469749, `RNS_PRIME_BITS'd566394243, `RNS_PRIME_BITS'd346619236, `RNS_PRIME_BITS'd448209918},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1348833947, `RNS_PRIME_BITS'd1844851629, `RNS_PRIME_BITS'd2004456777, `RNS_PRIME_BITS'd235031445, `RNS_PRIME_BITS'd1735102741, `RNS_PRIME_BITS'd583972638, `RNS_PRIME_BITS'd1580030603, `RNS_PRIME_BITS'd1054953566, `RNS_PRIME_BITS'd2062421468, `RNS_PRIME_BITS'd1048344043},
			'{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd1345114424, `RNS_PRIME_BITS'd1302007359, `RNS_PRIME_BITS'd92577089, `RNS_PRIME_BITS'd1971604877, `RNS_PRIME_BITS'd575557263, `RNS_PRIME_BITS'd2102231964, `RNS_PRIME_BITS'd967102215, `RNS_PRIME_BITS'd904263817, `RNS_PRIME_BITS'd592154024, `RNS_PRIME_BITS'd1495857983},
			'{`RNS_PRIME_BITS'd66, `RNS_PRIME_BITS'd637489359, `RNS_PRIME_BITS'd1479558466, `RNS_PRIME_BITS'd1903969447, `RNS_PRIME_BITS'd1183319220, `RNS_PRIME_BITS'd908246980, `RNS_PRIME_BITS'd1332127260, `RNS_PRIME_BITS'd11498795, `RNS_PRIME_BITS'd1231585878, `RNS_PRIME_BITS'd863775577, `RNS_PRIME_BITS'd1464649121},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd890668921, `RNS_PRIME_BITS'd1929701503, `RNS_PRIME_BITS'd1114795254, `RNS_PRIME_BITS'd1131199896, `RNS_PRIME_BITS'd1413802139, `RNS_PRIME_BITS'd1787419913, `RNS_PRIME_BITS'd285329909, `RNS_PRIME_BITS'd532056630, `RNS_PRIME_BITS'd1696529244, `RNS_PRIME_BITS'd1141319206},
			'{`RNS_PRIME_BITS'd254, `RNS_PRIME_BITS'd1628529615, `RNS_PRIME_BITS'd1072570713, `RNS_PRIME_BITS'd1400515486, `RNS_PRIME_BITS'd1033371745, `RNS_PRIME_BITS'd142818692, `RNS_PRIME_BITS'd635409143, `RNS_PRIME_BITS'd1555605954, `RNS_PRIME_BITS'd65591225, `RNS_PRIME_BITS'd51494655, `RNS_PRIME_BITS'd185332239},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd559630670, `RNS_PRIME_BITS'd269234662, `RNS_PRIME_BITS'd1139481071, `RNS_PRIME_BITS'd1776376047, `RNS_PRIME_BITS'd256922405, `RNS_PRIME_BITS'd352229326, `RNS_PRIME_BITS'd367110130, `RNS_PRIME_BITS'd2109514594, `RNS_PRIME_BITS'd452879539, `RNS_PRIME_BITS'd1521114358},
			'{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd1157501329, `RNS_PRIME_BITS'd1171055296, `RNS_PRIME_BITS'd243161416, `RNS_PRIME_BITS'd736480290, `RNS_PRIME_BITS'd546137976, `RNS_PRIME_BITS'd1040159993, `RNS_PRIME_BITS'd789556556, `RNS_PRIME_BITS'd1909978578, `RNS_PRIME_BITS'd899211686, `RNS_PRIME_BITS'd810246693},
			'{`RNS_PRIME_BITS'd220, `RNS_PRIME_BITS'd913953323, `RNS_PRIME_BITS'd166630647, `RNS_PRIME_BITS'd794861792, `RNS_PRIME_BITS'd1308251555, `RNS_PRIME_BITS'd220024834, `RNS_PRIME_BITS'd2067090424, `RNS_PRIME_BITS'd1895123462, `RNS_PRIME_BITS'd736098302, `RNS_PRIME_BITS'd1650113038, `RNS_PRIME_BITS'd1811599151},
			'{`RNS_PRIME_BITS'd230, `RNS_PRIME_BITS'd25314846, `RNS_PRIME_BITS'd1344453719, `RNS_PRIME_BITS'd1990288460, `RNS_PRIME_BITS'd1286263876, `RNS_PRIME_BITS'd1850587102, `RNS_PRIME_BITS'd726074958, `RNS_PRIME_BITS'd864152023, `RNS_PRIME_BITS'd120912832, `RNS_PRIME_BITS'd665760858, `RNS_PRIME_BITS'd2060756164},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1791644713, `RNS_PRIME_BITS'd161712777, `RNS_PRIME_BITS'd1295353801, `RNS_PRIME_BITS'd527998255, `RNS_PRIME_BITS'd508704, `RNS_PRIME_BITS'd1638712404, `RNS_PRIME_BITS'd887329497, `RNS_PRIME_BITS'd132166131, `RNS_PRIME_BITS'd624670822, `RNS_PRIME_BITS'd242506097},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd589099632, `RNS_PRIME_BITS'd1440836908, `RNS_PRIME_BITS'd1716054161, `RNS_PRIME_BITS'd1024915296, `RNS_PRIME_BITS'd334144567, `RNS_PRIME_BITS'd227492620, `RNS_PRIME_BITS'd1863095083, `RNS_PRIME_BITS'd845646242, `RNS_PRIME_BITS'd1809847005, `RNS_PRIME_BITS'd113316753},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd1339076758, `RNS_PRIME_BITS'd769734859, `RNS_PRIME_BITS'd1539848123, `RNS_PRIME_BITS'd1446728914, `RNS_PRIME_BITS'd747498299, `RNS_PRIME_BITS'd1395448515, `RNS_PRIME_BITS'd483453344, `RNS_PRIME_BITS'd107117875, `RNS_PRIME_BITS'd2064707598, `RNS_PRIME_BITS'd1091483909},
			'{`RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd1257537277, `RNS_PRIME_BITS'd1362879338, `RNS_PRIME_BITS'd940297036, `RNS_PRIME_BITS'd1572807336, `RNS_PRIME_BITS'd1479546086, `RNS_PRIME_BITS'd1951134535, `RNS_PRIME_BITS'd595248706, `RNS_PRIME_BITS'd654549710, `RNS_PRIME_BITS'd735033161, `RNS_PRIME_BITS'd1217965778},
			'{`RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd1114307253, `RNS_PRIME_BITS'd1065859291, `RNS_PRIME_BITS'd59885519, `RNS_PRIME_BITS'd690847805, `RNS_PRIME_BITS'd486609063, `RNS_PRIME_BITS'd1233411043, `RNS_PRIME_BITS'd955506154, `RNS_PRIME_BITS'd1013817448, `RNS_PRIME_BITS'd288658942, `RNS_PRIME_BITS'd1875894412},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd107566261, `RNS_PRIME_BITS'd535379015, `RNS_PRIME_BITS'd1349744976, `RNS_PRIME_BITS'd923272612, `RNS_PRIME_BITS'd241847474, `RNS_PRIME_BITS'd1194835589, `RNS_PRIME_BITS'd1822601058, `RNS_PRIME_BITS'd162506953, `RNS_PRIME_BITS'd1487954239, `RNS_PRIME_BITS'd172735353},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd152044712, `RNS_PRIME_BITS'd1717974170, `RNS_PRIME_BITS'd1177368815, `RNS_PRIME_BITS'd2032048140, `RNS_PRIME_BITS'd541265162, `RNS_PRIME_BITS'd2111205579, `RNS_PRIME_BITS'd1336457058, `RNS_PRIME_BITS'd275964119, `RNS_PRIME_BITS'd1185838874, `RNS_PRIME_BITS'd971052263},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd923748325, `RNS_PRIME_BITS'd1359015913, `RNS_PRIME_BITS'd1370508929, `RNS_PRIME_BITS'd1073464063, `RNS_PRIME_BITS'd1626464979, `RNS_PRIME_BITS'd62055301, `RNS_PRIME_BITS'd35341169, `RNS_PRIME_BITS'd648759873, `RNS_PRIME_BITS'd1627653868, `RNS_PRIME_BITS'd1633532570},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd1968764293, `RNS_PRIME_BITS'd625254340, `RNS_PRIME_BITS'd1928932687, `RNS_PRIME_BITS'd263818109, `RNS_PRIME_BITS'd1403738007, `RNS_PRIME_BITS'd1715138468, `RNS_PRIME_BITS'd994309017, `RNS_PRIME_BITS'd326940506, `RNS_PRIME_BITS'd2044618763, `RNS_PRIME_BITS'd853289331},
			'{`RNS_PRIME_BITS'd189, `RNS_PRIME_BITS'd723421897, `RNS_PRIME_BITS'd1080926945, `RNS_PRIME_BITS'd1140924078, `RNS_PRIME_BITS'd223602630, `RNS_PRIME_BITS'd1292075945, `RNS_PRIME_BITS'd1289017984, `RNS_PRIME_BITS'd1769819368, `RNS_PRIME_BITS'd1326090145, `RNS_PRIME_BITS'd1845654709, `RNS_PRIME_BITS'd838360829},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd1519989365, `RNS_PRIME_BITS'd65234468, `RNS_PRIME_BITS'd972169002, `RNS_PRIME_BITS'd814267858, `RNS_PRIME_BITS'd3501337, `RNS_PRIME_BITS'd1805339177, `RNS_PRIME_BITS'd118876390, `RNS_PRIME_BITS'd1335138655, `RNS_PRIME_BITS'd2033426768, `RNS_PRIME_BITS'd2142951653},
			'{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd15650524, `RNS_PRIME_BITS'd1293822637, `RNS_PRIME_BITS'd1662710961, `RNS_PRIME_BITS'd1744198421, `RNS_PRIME_BITS'd760925998, `RNS_PRIME_BITS'd1990310669, `RNS_PRIME_BITS'd720457635, `RNS_PRIME_BITS'd879535769, `RNS_PRIME_BITS'd1109288995, `RNS_PRIME_BITS'd1098886785},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd802459139, `RNS_PRIME_BITS'd1862062953, `RNS_PRIME_BITS'd951545330, `RNS_PRIME_BITS'd860848899, `RNS_PRIME_BITS'd1079246348, `RNS_PRIME_BITS'd1537499607, `RNS_PRIME_BITS'd1336360573, `RNS_PRIME_BITS'd1558253840, `RNS_PRIME_BITS'd525161866, `RNS_PRIME_BITS'd1730630972},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd306569084, `RNS_PRIME_BITS'd1840021757, `RNS_PRIME_BITS'd1640478532, `RNS_PRIME_BITS'd1301738641, `RNS_PRIME_BITS'd266624620, `RNS_PRIME_BITS'd1587949734, `RNS_PRIME_BITS'd1677462924, `RNS_PRIME_BITS'd1102874180, `RNS_PRIME_BITS'd2044943950, `RNS_PRIME_BITS'd690302665},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd233370496, `RNS_PRIME_BITS'd1800291942, `RNS_PRIME_BITS'd682154649, `RNS_PRIME_BITS'd1368041010, `RNS_PRIME_BITS'd791285229, `RNS_PRIME_BITS'd1289022131, `RNS_PRIME_BITS'd1406320158, `RNS_PRIME_BITS'd1557631444, `RNS_PRIME_BITS'd32834913, `RNS_PRIME_BITS'd902282165},
			'{`RNS_PRIME_BITS'd244, `RNS_PRIME_BITS'd240223384, `RNS_PRIME_BITS'd891844296, `RNS_PRIME_BITS'd1648909567, `RNS_PRIME_BITS'd1910006597, `RNS_PRIME_BITS'd259729073, `RNS_PRIME_BITS'd2125212460, `RNS_PRIME_BITS'd319171641, `RNS_PRIME_BITS'd597661704, `RNS_PRIME_BITS'd1331472727, `RNS_PRIME_BITS'd466572194},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd602783278, `RNS_PRIME_BITS'd306212216, `RNS_PRIME_BITS'd2024751924, `RNS_PRIME_BITS'd788173821, `RNS_PRIME_BITS'd401110859, `RNS_PRIME_BITS'd896568438, `RNS_PRIME_BITS'd1195528387, `RNS_PRIME_BITS'd1325317927, `RNS_PRIME_BITS'd1759550114, `RNS_PRIME_BITS'd1174991516},
			'{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd1506902842, `RNS_PRIME_BITS'd835139412, `RNS_PRIME_BITS'd1899202744, `RNS_PRIME_BITS'd578424927, `RNS_PRIME_BITS'd78737645, `RNS_PRIME_BITS'd1810375274, `RNS_PRIME_BITS'd1019945138, `RNS_PRIME_BITS'd1476494174, `RNS_PRIME_BITS'd1948825999, `RNS_PRIME_BITS'd1816413912},
			'{`RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd1955957184, `RNS_PRIME_BITS'd724421342, `RNS_PRIME_BITS'd778583987, `RNS_PRIME_BITS'd1504218104, `RNS_PRIME_BITS'd2136016041, `RNS_PRIME_BITS'd934268666, `RNS_PRIME_BITS'd1821958871, `RNS_PRIME_BITS'd656249630, `RNS_PRIME_BITS'd606860525, `RNS_PRIME_BITS'd1108050209},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd142480780, `RNS_PRIME_BITS'd1076951153, `RNS_PRIME_BITS'd1469737589, `RNS_PRIME_BITS'd888050255, `RNS_PRIME_BITS'd1138977787, `RNS_PRIME_BITS'd322674830, `RNS_PRIME_BITS'd715245453, `RNS_PRIME_BITS'd1082053094, `RNS_PRIME_BITS'd227722567, `RNS_PRIME_BITS'd1529541656},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1083236422, `RNS_PRIME_BITS'd1629772037, `RNS_PRIME_BITS'd421185093, `RNS_PRIME_BITS'd277875174, `RNS_PRIME_BITS'd836725873, `RNS_PRIME_BITS'd111119244, `RNS_PRIME_BITS'd1466670951, `RNS_PRIME_BITS'd1678899526, `RNS_PRIME_BITS'd332703821, `RNS_PRIME_BITS'd926564010},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1309966671, `RNS_PRIME_BITS'd958613410, `RNS_PRIME_BITS'd501501938, `RNS_PRIME_BITS'd532199149, `RNS_PRIME_BITS'd692929505, `RNS_PRIME_BITS'd837613327, `RNS_PRIME_BITS'd1414219209, `RNS_PRIME_BITS'd1998672519, `RNS_PRIME_BITS'd646058240, `RNS_PRIME_BITS'd376122387},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd1836229569, `RNS_PRIME_BITS'd795580179, `RNS_PRIME_BITS'd699906758, `RNS_PRIME_BITS'd1321942828, `RNS_PRIME_BITS'd1175498707, `RNS_PRIME_BITS'd1341561911, `RNS_PRIME_BITS'd3694551, `RNS_PRIME_BITS'd524241530, `RNS_PRIME_BITS'd870597670, `RNS_PRIME_BITS'd1255036559},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1820523574, `RNS_PRIME_BITS'd1209558314, `RNS_PRIME_BITS'd1191885383, `RNS_PRIME_BITS'd1099754634, `RNS_PRIME_BITS'd328855164, `RNS_PRIME_BITS'd397815075, `RNS_PRIME_BITS'd1704622002, `RNS_PRIME_BITS'd191375772, `RNS_PRIME_BITS'd637045312, `RNS_PRIME_BITS'd4148703},
			'{`RNS_PRIME_BITS'd76, `RNS_PRIME_BITS'd327232664, `RNS_PRIME_BITS'd400426857, `RNS_PRIME_BITS'd1599444619, `RNS_PRIME_BITS'd749735936, `RNS_PRIME_BITS'd1678896958, `RNS_PRIME_BITS'd1283180472, `RNS_PRIME_BITS'd1281999832, `RNS_PRIME_BITS'd1833558253, `RNS_PRIME_BITS'd707354233, `RNS_PRIME_BITS'd1948380049},
			'{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd2049882085, `RNS_PRIME_BITS'd2105210570, `RNS_PRIME_BITS'd12448303, `RNS_PRIME_BITS'd881555272, `RNS_PRIME_BITS'd1762730962, `RNS_PRIME_BITS'd1744916055, `RNS_PRIME_BITS'd794724046, `RNS_PRIME_BITS'd166030696, `RNS_PRIME_BITS'd482240971, `RNS_PRIME_BITS'd1000819526},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd354361265, `RNS_PRIME_BITS'd1494498431, `RNS_PRIME_BITS'd1919837893, `RNS_PRIME_BITS'd1107392755, `RNS_PRIME_BITS'd961102314, `RNS_PRIME_BITS'd1941116829, `RNS_PRIME_BITS'd1581130677, `RNS_PRIME_BITS'd2033788341, `RNS_PRIME_BITS'd1279223657, `RNS_PRIME_BITS'd441782404},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd1271901409, `RNS_PRIME_BITS'd138914877, `RNS_PRIME_BITS'd275616970, `RNS_PRIME_BITS'd1646120547, `RNS_PRIME_BITS'd115918287, `RNS_PRIME_BITS'd661140201, `RNS_PRIME_BITS'd1978364965, `RNS_PRIME_BITS'd1017107895, `RNS_PRIME_BITS'd1297149731, `RNS_PRIME_BITS'd1249075327},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1381289890, `RNS_PRIME_BITS'd2018184917, `RNS_PRIME_BITS'd902583850, `RNS_PRIME_BITS'd1700172634, `RNS_PRIME_BITS'd625015279, `RNS_PRIME_BITS'd628896427, `RNS_PRIME_BITS'd1444165050, `RNS_PRIME_BITS'd871763951, `RNS_PRIME_BITS'd117677784, `RNS_PRIME_BITS'd777001115},
			'{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd1246195080, `RNS_PRIME_BITS'd662445337, `RNS_PRIME_BITS'd420747815, `RNS_PRIME_BITS'd1075863020, `RNS_PRIME_BITS'd544827408, `RNS_PRIME_BITS'd1680249467, `RNS_PRIME_BITS'd1531537342, `RNS_PRIME_BITS'd901034090, `RNS_PRIME_BITS'd153316553, `RNS_PRIME_BITS'd1656237532},
			'{`RNS_PRIME_BITS'd69, `RNS_PRIME_BITS'd1647999649, `RNS_PRIME_BITS'd1771190978, `RNS_PRIME_BITS'd1694548415, `RNS_PRIME_BITS'd1840556195, `RNS_PRIME_BITS'd830534578, `RNS_PRIME_BITS'd1799590543, `RNS_PRIME_BITS'd1095917823, `RNS_PRIME_BITS'd2124984111, `RNS_PRIME_BITS'd76315630, `RNS_PRIME_BITS'd2114738654},
			'{`RNS_PRIME_BITS'd14, `RNS_PRIME_BITS'd1291008316, `RNS_PRIME_BITS'd1510124479, `RNS_PRIME_BITS'd697967636, `RNS_PRIME_BITS'd1683137498, `RNS_PRIME_BITS'd512431576, `RNS_PRIME_BITS'd510160379, `RNS_PRIME_BITS'd1383153078, `RNS_PRIME_BITS'd1091355969, `RNS_PRIME_BITS'd1516202209, `RNS_PRIME_BITS'd1719247936},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd1201016571, `RNS_PRIME_BITS'd528807111, `RNS_PRIME_BITS'd1876010778, `RNS_PRIME_BITS'd1042483073, `RNS_PRIME_BITS'd1238318331, `RNS_PRIME_BITS'd1382860398, `RNS_PRIME_BITS'd1757241977, `RNS_PRIME_BITS'd912580083, `RNS_PRIME_BITS'd1527393628, `RNS_PRIME_BITS'd350941306},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd1421615102, `RNS_PRIME_BITS'd284313799, `RNS_PRIME_BITS'd1742428325, `RNS_PRIME_BITS'd1686394895, `RNS_PRIME_BITS'd1615779245, `RNS_PRIME_BITS'd319208443, `RNS_PRIME_BITS'd1525115317, `RNS_PRIME_BITS'd592536841, `RNS_PRIME_BITS'd932528472, `RNS_PRIME_BITS'd1551338288},
			'{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd17637367, `RNS_PRIME_BITS'd1562399507, `RNS_PRIME_BITS'd1435510522, `RNS_PRIME_BITS'd469108704, `RNS_PRIME_BITS'd542199375, `RNS_PRIME_BITS'd918147342, `RNS_PRIME_BITS'd149614217, `RNS_PRIME_BITS'd2141828327, `RNS_PRIME_BITS'd1883145958, `RNS_PRIME_BITS'd300987089},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd1157734352, `RNS_PRIME_BITS'd1854124505, `RNS_PRIME_BITS'd513731701, `RNS_PRIME_BITS'd1682857761, `RNS_PRIME_BITS'd334414650, `RNS_PRIME_BITS'd953965897, `RNS_PRIME_BITS'd1006718855, `RNS_PRIME_BITS'd532530418, `RNS_PRIME_BITS'd815315064, `RNS_PRIME_BITS'd1969632419},
			'{`RNS_PRIME_BITS'd40, `RNS_PRIME_BITS'd2117482484, `RNS_PRIME_BITS'd2061709753, `RNS_PRIME_BITS'd518509583, `RNS_PRIME_BITS'd2097930504, `RNS_PRIME_BITS'd2144922307, `RNS_PRIME_BITS'd131968939, `RNS_PRIME_BITS'd1347107026, `RNS_PRIME_BITS'd77762930, `RNS_PRIME_BITS'd1440623138, `RNS_PRIME_BITS'd1172492088},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd1816686281, `RNS_PRIME_BITS'd866875819, `RNS_PRIME_BITS'd591543259, `RNS_PRIME_BITS'd2086870251, `RNS_PRIME_BITS'd1600950822, `RNS_PRIME_BITS'd2110102715, `RNS_PRIME_BITS'd117299070, `RNS_PRIME_BITS'd577232477, `RNS_PRIME_BITS'd257154307, `RNS_PRIME_BITS'd1441407288},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd1158338557, `RNS_PRIME_BITS'd159455344, `RNS_PRIME_BITS'd1640935915, `RNS_PRIME_BITS'd1075683447, `RNS_PRIME_BITS'd1642852325, `RNS_PRIME_BITS'd73123535, `RNS_PRIME_BITS'd1918977663, `RNS_PRIME_BITS'd2031710906, `RNS_PRIME_BITS'd464398154, `RNS_PRIME_BITS'd2044522004},
			'{`RNS_PRIME_BITS'd200, `RNS_PRIME_BITS'd697831407, `RNS_PRIME_BITS'd286548012, `RNS_PRIME_BITS'd1973402441, `RNS_PRIME_BITS'd97280642, `RNS_PRIME_BITS'd959862771, `RNS_PRIME_BITS'd2107610452, `RNS_PRIME_BITS'd1273143702, `RNS_PRIME_BITS'd875705394, `RNS_PRIME_BITS'd1656305303, `RNS_PRIME_BITS'd890105596},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd1249949978, `RNS_PRIME_BITS'd1571138432, `RNS_PRIME_BITS'd1720591807, `RNS_PRIME_BITS'd170538012, `RNS_PRIME_BITS'd139069934, `RNS_PRIME_BITS'd2124247611, `RNS_PRIME_BITS'd128204835, `RNS_PRIME_BITS'd67401812, `RNS_PRIME_BITS'd149186395, `RNS_PRIME_BITS'd981922731},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd707035355, `RNS_PRIME_BITS'd1600460038, `RNS_PRIME_BITS'd884764309, `RNS_PRIME_BITS'd1489459444, `RNS_PRIME_BITS'd1053381919, `RNS_PRIME_BITS'd677138648, `RNS_PRIME_BITS'd1560660816, `RNS_PRIME_BITS'd1796904162, `RNS_PRIME_BITS'd1070114158, `RNS_PRIME_BITS'd1711156906},
			'{`RNS_PRIME_BITS'd127, `RNS_PRIME_BITS'd1621024850, `RNS_PRIME_BITS'd968139671, `RNS_PRIME_BITS'd161554646, `RNS_PRIME_BITS'd1435692300, `RNS_PRIME_BITS'd479351687, `RNS_PRIME_BITS'd1267909006, `RNS_PRIME_BITS'd555104894, `RNS_PRIME_BITS'd379659211, `RNS_PRIME_BITS'd714606488, `RNS_PRIME_BITS'd1145928960},
			'{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd306271144, `RNS_PRIME_BITS'd1768009783, `RNS_PRIME_BITS'd2009184009, `RNS_PRIME_BITS'd2141804236, `RNS_PRIME_BITS'd1641508139, `RNS_PRIME_BITS'd1960129629, `RNS_PRIME_BITS'd646433138, `RNS_PRIME_BITS'd81594901, `RNS_PRIME_BITS'd265317, `RNS_PRIME_BITS'd1611337738},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd258113990, `RNS_PRIME_BITS'd2039434436, `RNS_PRIME_BITS'd1261611557, `RNS_PRIME_BITS'd1780956481, `RNS_PRIME_BITS'd1463875624, `RNS_PRIME_BITS'd1349684416, `RNS_PRIME_BITS'd1888810822, `RNS_PRIME_BITS'd1652095714, `RNS_PRIME_BITS'd1255250998, `RNS_PRIME_BITS'd775078885},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd1221198069, `RNS_PRIME_BITS'd2143116151, `RNS_PRIME_BITS'd1592556941, `RNS_PRIME_BITS'd34435693, `RNS_PRIME_BITS'd1533194705, `RNS_PRIME_BITS'd394551915, `RNS_PRIME_BITS'd1285881103, `RNS_PRIME_BITS'd470486345, `RNS_PRIME_BITS'd622453981, `RNS_PRIME_BITS'd627239343},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd618098919, `RNS_PRIME_BITS'd238087225, `RNS_PRIME_BITS'd447382298, `RNS_PRIME_BITS'd352302497, `RNS_PRIME_BITS'd1996607689, `RNS_PRIME_BITS'd913606149, `RNS_PRIME_BITS'd1850984129, `RNS_PRIME_BITS'd342824710, `RNS_PRIME_BITS'd1390425313, `RNS_PRIME_BITS'd1430369291},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd423200828, `RNS_PRIME_BITS'd1648540232, `RNS_PRIME_BITS'd992856097, `RNS_PRIME_BITS'd2058280730, `RNS_PRIME_BITS'd129063228, `RNS_PRIME_BITS'd1015186439, `RNS_PRIME_BITS'd1012379207, `RNS_PRIME_BITS'd343789635, `RNS_PRIME_BITS'd331955084, `RNS_PRIME_BITS'd917353169},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd1850589253, `RNS_PRIME_BITS'd1621717790, `RNS_PRIME_BITS'd541920963, `RNS_PRIME_BITS'd1809565732, `RNS_PRIME_BITS'd1183718773, `RNS_PRIME_BITS'd686718554, `RNS_PRIME_BITS'd1676366113, `RNS_PRIME_BITS'd117706650, `RNS_PRIME_BITS'd1418630883, `RNS_PRIME_BITS'd1539299055},
			'{`RNS_PRIME_BITS'd152, `RNS_PRIME_BITS'd401963463, `RNS_PRIME_BITS'd1015901580, `RNS_PRIME_BITS'd850298754, `RNS_PRIME_BITS'd1612974951, `RNS_PRIME_BITS'd1245244323, `RNS_PRIME_BITS'd1539882473, `RNS_PRIME_BITS'd770310686, `RNS_PRIME_BITS'd532798600, `RNS_PRIME_BITS'd762020549, `RNS_PRIME_BITS'd364826689}
		},
		'{
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd496664282, `RNS_PRIME_BITS'd1363778345, `RNS_PRIME_BITS'd1035556982, `RNS_PRIME_BITS'd805578265, `RNS_PRIME_BITS'd549166752, `RNS_PRIME_BITS'd1574666888, `RNS_PRIME_BITS'd1858496281, `RNS_PRIME_BITS'd1007870612, `RNS_PRIME_BITS'd227114546, `RNS_PRIME_BITS'd1793606260},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1608567105, `RNS_PRIME_BITS'd1529058673, `RNS_PRIME_BITS'd808973517, `RNS_PRIME_BITS'd130845307, `RNS_PRIME_BITS'd50117541, `RNS_PRIME_BITS'd122361920, `RNS_PRIME_BITS'd596466224, `RNS_PRIME_BITS'd1107797424, `RNS_PRIME_BITS'd185656935, `RNS_PRIME_BITS'd789787990},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1337484787, `RNS_PRIME_BITS'd57962201, `RNS_PRIME_BITS'd546299570, `RNS_PRIME_BITS'd1300802353, `RNS_PRIME_BITS'd204518873, `RNS_PRIME_BITS'd1242686070, `RNS_PRIME_BITS'd618756376, `RNS_PRIME_BITS'd1460113389, `RNS_PRIME_BITS'd2096650530, `RNS_PRIME_BITS'd859568432},
			'{`RNS_PRIME_BITS'd40, `RNS_PRIME_BITS'd444205039, `RNS_PRIME_BITS'd1628533368, `RNS_PRIME_BITS'd1782321273, `RNS_PRIME_BITS'd971211237, `RNS_PRIME_BITS'd1549754476, `RNS_PRIME_BITS'd1841296949, `RNS_PRIME_BITS'd686579453, `RNS_PRIME_BITS'd331572205, `RNS_PRIME_BITS'd329692279, `RNS_PRIME_BITS'd462204125},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1445398008, `RNS_PRIME_BITS'd653456047, `RNS_PRIME_BITS'd35482018, `RNS_PRIME_BITS'd557496536, `RNS_PRIME_BITS'd267790300, `RNS_PRIME_BITS'd843176199, `RNS_PRIME_BITS'd227928720, `RNS_PRIME_BITS'd1264273532, `RNS_PRIME_BITS'd235239605, `RNS_PRIME_BITS'd771311141},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd1666181169, `RNS_PRIME_BITS'd160514543, `RNS_PRIME_BITS'd1399676730, `RNS_PRIME_BITS'd1097639396, `RNS_PRIME_BITS'd942268911, `RNS_PRIME_BITS'd1088925803, `RNS_PRIME_BITS'd2144239244, `RNS_PRIME_BITS'd924622711, `RNS_PRIME_BITS'd270820994, `RNS_PRIME_BITS'd110273218},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd1244971827, `RNS_PRIME_BITS'd46221564, `RNS_PRIME_BITS'd262500625, `RNS_PRIME_BITS'd639584943, `RNS_PRIME_BITS'd306540021, `RNS_PRIME_BITS'd1912552501, `RNS_PRIME_BITS'd1073679567, `RNS_PRIME_BITS'd713904558, `RNS_PRIME_BITS'd268372791, `RNS_PRIME_BITS'd191841818},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd698318862, `RNS_PRIME_BITS'd232734665, `RNS_PRIME_BITS'd192363136, `RNS_PRIME_BITS'd488675673, `RNS_PRIME_BITS'd1981601082, `RNS_PRIME_BITS'd1213634479, `RNS_PRIME_BITS'd647079262, `RNS_PRIME_BITS'd1067173597, `RNS_PRIME_BITS'd641660871, `RNS_PRIME_BITS'd1921190254},
			'{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd2066114937, `RNS_PRIME_BITS'd1459847815, `RNS_PRIME_BITS'd1289319664, `RNS_PRIME_BITS'd1804854032, `RNS_PRIME_BITS'd111944773, `RNS_PRIME_BITS'd2097774118, `RNS_PRIME_BITS'd100423507, `RNS_PRIME_BITS'd91312048, `RNS_PRIME_BITS'd2114801649, `RNS_PRIME_BITS'd18894692},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1914187354, `RNS_PRIME_BITS'd1774684653, `RNS_PRIME_BITS'd1513894601, `RNS_PRIME_BITS'd925092001, `RNS_PRIME_BITS'd1061825663, `RNS_PRIME_BITS'd1754979706, `RNS_PRIME_BITS'd2120919600, `RNS_PRIME_BITS'd1728507285, `RNS_PRIME_BITS'd835252734, `RNS_PRIME_BITS'd1036996988},
			'{`RNS_PRIME_BITS'd160, `RNS_PRIME_BITS'd392076842, `RNS_PRIME_BITS'd908438224, `RNS_PRIME_BITS'd861154708, `RNS_PRIME_BITS'd1107818706, `RNS_PRIME_BITS'd256742250, `RNS_PRIME_BITS'd895682518, `RNS_PRIME_BITS'd389732213, `RNS_PRIME_BITS'd929274275, `RNS_PRIME_BITS'd513243327, `RNS_PRIME_BITS'd924769361},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd651434042, `RNS_PRIME_BITS'd584858919, `RNS_PRIME_BITS'd1568165086, `RNS_PRIME_BITS'd135842525, `RNS_PRIME_BITS'd200347940, `RNS_PRIME_BITS'd927071129, `RNS_PRIME_BITS'd422159745, `RNS_PRIME_BITS'd1076108391, `RNS_PRIME_BITS'd77951812, `RNS_PRIME_BITS'd145555725},
			'{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd715951950, `RNS_PRIME_BITS'd1914156239, `RNS_PRIME_BITS'd1135832849, `RNS_PRIME_BITS'd447445819, `RNS_PRIME_BITS'd1768578018, `RNS_PRIME_BITS'd1755827369, `RNS_PRIME_BITS'd59844739, `RNS_PRIME_BITS'd1166576027, `RNS_PRIME_BITS'd1223204782, `RNS_PRIME_BITS'd1795161428},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd1937925685, `RNS_PRIME_BITS'd636733489, `RNS_PRIME_BITS'd1093154378, `RNS_PRIME_BITS'd646090295, `RNS_PRIME_BITS'd2095744800, `RNS_PRIME_BITS'd1235273673, `RNS_PRIME_BITS'd1939374608, `RNS_PRIME_BITS'd1232318059, `RNS_PRIME_BITS'd2056395400, `RNS_PRIME_BITS'd542063678},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd592528257, `RNS_PRIME_BITS'd4554121, `RNS_PRIME_BITS'd752596956, `RNS_PRIME_BITS'd1999520000, `RNS_PRIME_BITS'd1735588202, `RNS_PRIME_BITS'd486970230, `RNS_PRIME_BITS'd1609555766, `RNS_PRIME_BITS'd2050423213, `RNS_PRIME_BITS'd1636767231, `RNS_PRIME_BITS'd1372805036},
			'{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd1890304033, `RNS_PRIME_BITS'd1626537980, `RNS_PRIME_BITS'd1535419953, `RNS_PRIME_BITS'd1914748354, `RNS_PRIME_BITS'd858438522, `RNS_PRIME_BITS'd97096333, `RNS_PRIME_BITS'd1143059163, `RNS_PRIME_BITS'd684949220, `RNS_PRIME_BITS'd1437767108, `RNS_PRIME_BITS'd1838378478},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd160721397, `RNS_PRIME_BITS'd1165722807, `RNS_PRIME_BITS'd178613915, `RNS_PRIME_BITS'd618542610, `RNS_PRIME_BITS'd1737671766, `RNS_PRIME_BITS'd1249208216, `RNS_PRIME_BITS'd546719219, `RNS_PRIME_BITS'd1955667676, `RNS_PRIME_BITS'd2137285411, `RNS_PRIME_BITS'd418147965},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd1692665063, `RNS_PRIME_BITS'd33890232, `RNS_PRIME_BITS'd1009185866, `RNS_PRIME_BITS'd1536228269, `RNS_PRIME_BITS'd1852054839, `RNS_PRIME_BITS'd326639357, `RNS_PRIME_BITS'd49948394, `RNS_PRIME_BITS'd1775330783, `RNS_PRIME_BITS'd341529866, `RNS_PRIME_BITS'd1416326890},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd546941176, `RNS_PRIME_BITS'd1243326244, `RNS_PRIME_BITS'd556627411, `RNS_PRIME_BITS'd748055092, `RNS_PRIME_BITS'd249328861, `RNS_PRIME_BITS'd645331390, `RNS_PRIME_BITS'd1378628194, `RNS_PRIME_BITS'd1351865321, `RNS_PRIME_BITS'd76682022, `RNS_PRIME_BITS'd1192143176},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd130004873, `RNS_PRIME_BITS'd2044909686, `RNS_PRIME_BITS'd2056059945, `RNS_PRIME_BITS'd1641827291, `RNS_PRIME_BITS'd645928843, `RNS_PRIME_BITS'd940067925, `RNS_PRIME_BITS'd1626038, `RNS_PRIME_BITS'd67558171, `RNS_PRIME_BITS'd1177336351, `RNS_PRIME_BITS'd1030798525},
			'{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd789957968, `RNS_PRIME_BITS'd487554740, `RNS_PRIME_BITS'd1818409103, `RNS_PRIME_BITS'd1742687747, `RNS_PRIME_BITS'd1228414497, `RNS_PRIME_BITS'd1356870324, `RNS_PRIME_BITS'd1403700268, `RNS_PRIME_BITS'd172255780, `RNS_PRIME_BITS'd492317479, `RNS_PRIME_BITS'd451057652},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd715064509, `RNS_PRIME_BITS'd228761151, `RNS_PRIME_BITS'd2000507384, `RNS_PRIME_BITS'd1536858362, `RNS_PRIME_BITS'd1433758064, `RNS_PRIME_BITS'd1225416533, `RNS_PRIME_BITS'd627282315, `RNS_PRIME_BITS'd2105694895, `RNS_PRIME_BITS'd143108326, `RNS_PRIME_BITS'd1103218755},
			'{`RNS_PRIME_BITS'd12, `RNS_PRIME_BITS'd1005291939, `RNS_PRIME_BITS'd1129282534, `RNS_PRIME_BITS'd1948622800, `RNS_PRIME_BITS'd95687708, `RNS_PRIME_BITS'd1546513386, `RNS_PRIME_BITS'd2036072794, `RNS_PRIME_BITS'd196371900, `RNS_PRIME_BITS'd1470580662, `RNS_PRIME_BITS'd616006809, `RNS_PRIME_BITS'd299036250},
			'{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd1980210264, `RNS_PRIME_BITS'd1834024258, `RNS_PRIME_BITS'd877384359, `RNS_PRIME_BITS'd1106481895, `RNS_PRIME_BITS'd1540005035, `RNS_PRIME_BITS'd1277135415, `RNS_PRIME_BITS'd822531474, `RNS_PRIME_BITS'd1256934628, `RNS_PRIME_BITS'd464248368, `RNS_PRIME_BITS'd1772677581},
			'{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd1130619139, `RNS_PRIME_BITS'd1097979843, `RNS_PRIME_BITS'd604560359, `RNS_PRIME_BITS'd212231565, `RNS_PRIME_BITS'd574977836, `RNS_PRIME_BITS'd1871836745, `RNS_PRIME_BITS'd1254861632, `RNS_PRIME_BITS'd162561079, `RNS_PRIME_BITS'd1658125439, `RNS_PRIME_BITS'd1509790644},
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd273214037, `RNS_PRIME_BITS'd2069372070, `RNS_PRIME_BITS'd1256531473, `RNS_PRIME_BITS'd1428753586, `RNS_PRIME_BITS'd49173564, `RNS_PRIME_BITS'd1075852553, `RNS_PRIME_BITS'd250170744, `RNS_PRIME_BITS'd309596760, `RNS_PRIME_BITS'd736634378, `RNS_PRIME_BITS'd224074578},
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd1541478806, `RNS_PRIME_BITS'd702345230, `RNS_PRIME_BITS'd283449234, `RNS_PRIME_BITS'd380257656, `RNS_PRIME_BITS'd594474276, `RNS_PRIME_BITS'd1910069111, `RNS_PRIME_BITS'd1807428007, `RNS_PRIME_BITS'd960962972, `RNS_PRIME_BITS'd1443695735, `RNS_PRIME_BITS'd1779472081},
			'{`RNS_PRIME_BITS'd12, `RNS_PRIME_BITS'd137429434, `RNS_PRIME_BITS'd457069847, `RNS_PRIME_BITS'd1208432458, `RNS_PRIME_BITS'd428123300, `RNS_PRIME_BITS'd1620499274, `RNS_PRIME_BITS'd2135310823, `RNS_PRIME_BITS'd384770328, `RNS_PRIME_BITS'd478679174, `RNS_PRIME_BITS'd1157247986, `RNS_PRIME_BITS'd1582187797},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd570612190, `RNS_PRIME_BITS'd1799770100, `RNS_PRIME_BITS'd1030378198, `RNS_PRIME_BITS'd2122628974, `RNS_PRIME_BITS'd1634202550, `RNS_PRIME_BITS'd100939365, `RNS_PRIME_BITS'd2067835945, `RNS_PRIME_BITS'd709725221, `RNS_PRIME_BITS'd425607033, `RNS_PRIME_BITS'd1274142585},
			'{`RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd338657896, `RNS_PRIME_BITS'd783358596, `RNS_PRIME_BITS'd2068335702, `RNS_PRIME_BITS'd556837996, `RNS_PRIME_BITS'd616302645, `RNS_PRIME_BITS'd529312369, `RNS_PRIME_BITS'd1457701368, `RNS_PRIME_BITS'd231985731, `RNS_PRIME_BITS'd3482439, `RNS_PRIME_BITS'd1016573947},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1416754925, `RNS_PRIME_BITS'd1545733734, `RNS_PRIME_BITS'd1341543566, `RNS_PRIME_BITS'd1292838522, `RNS_PRIME_BITS'd1189324473, `RNS_PRIME_BITS'd1370164736, `RNS_PRIME_BITS'd1947434612, `RNS_PRIME_BITS'd1086476724, `RNS_PRIME_BITS'd2085797309, `RNS_PRIME_BITS'd1166407585},
			'{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd269003453, `RNS_PRIME_BITS'd1620713953, `RNS_PRIME_BITS'd834067416, `RNS_PRIME_BITS'd1052904626, `RNS_PRIME_BITS'd866608925, `RNS_PRIME_BITS'd1832314288, `RNS_PRIME_BITS'd70423472, `RNS_PRIME_BITS'd1350498046, `RNS_PRIME_BITS'd1185610035, `RNS_PRIME_BITS'd29407452},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd1224156218, `RNS_PRIME_BITS'd737051057, `RNS_PRIME_BITS'd318215709, `RNS_PRIME_BITS'd701128438, `RNS_PRIME_BITS'd77872242, `RNS_PRIME_BITS'd1748197658, `RNS_PRIME_BITS'd599971828, `RNS_PRIME_BITS'd408942692, `RNS_PRIME_BITS'd1964881296, `RNS_PRIME_BITS'd1413509834},
			'{`RNS_PRIME_BITS'd220, `RNS_PRIME_BITS'd473450255, `RNS_PRIME_BITS'd78139058, `RNS_PRIME_BITS'd1781249803, `RNS_PRIME_BITS'd616335536, `RNS_PRIME_BITS'd1985723146, `RNS_PRIME_BITS'd989929804, `RNS_PRIME_BITS'd339804399, `RNS_PRIME_BITS'd1266133662, `RNS_PRIME_BITS'd1303938637, `RNS_PRIME_BITS'd378243656},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1703680388, `RNS_PRIME_BITS'd1990555555, `RNS_PRIME_BITS'd1598929657, `RNS_PRIME_BITS'd1821369459, `RNS_PRIME_BITS'd2030084534, `RNS_PRIME_BITS'd1532559916, `RNS_PRIME_BITS'd1763039863, `RNS_PRIME_BITS'd625230523, `RNS_PRIME_BITS'd964439729, `RNS_PRIME_BITS'd538831998},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd424603248, `RNS_PRIME_BITS'd1579373321, `RNS_PRIME_BITS'd361344986, `RNS_PRIME_BITS'd1465918973, `RNS_PRIME_BITS'd1965712374, `RNS_PRIME_BITS'd1745555260, `RNS_PRIME_BITS'd1203578436, `RNS_PRIME_BITS'd501049973, `RNS_PRIME_BITS'd1584558739, `RNS_PRIME_BITS'd2090336497},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1491492881, `RNS_PRIME_BITS'd2083048416, `RNS_PRIME_BITS'd1029662195, `RNS_PRIME_BITS'd1946096068, `RNS_PRIME_BITS'd1333004056, `RNS_PRIME_BITS'd270095625, `RNS_PRIME_BITS'd325578655, `RNS_PRIME_BITS'd1865616522, `RNS_PRIME_BITS'd1374309910, `RNS_PRIME_BITS'd1397456179},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd1305567534, `RNS_PRIME_BITS'd413125765, `RNS_PRIME_BITS'd810059952, `RNS_PRIME_BITS'd1456250738, `RNS_PRIME_BITS'd1386805384, `RNS_PRIME_BITS'd383613919, `RNS_PRIME_BITS'd252081990, `RNS_PRIME_BITS'd406541223, `RNS_PRIME_BITS'd1165791535, `RNS_PRIME_BITS'd876180326},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd763994593, `RNS_PRIME_BITS'd1310985626, `RNS_PRIME_BITS'd1806568640, `RNS_PRIME_BITS'd489820213, `RNS_PRIME_BITS'd2105285801, `RNS_PRIME_BITS'd1086946486, `RNS_PRIME_BITS'd1774486735, `RNS_PRIME_BITS'd1732766984, `RNS_PRIME_BITS'd241796333, `RNS_PRIME_BITS'd376420771},
			'{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd105842390, `RNS_PRIME_BITS'd1556655645, `RNS_PRIME_BITS'd1640859800, `RNS_PRIME_BITS'd895436980, `RNS_PRIME_BITS'd2146580905, `RNS_PRIME_BITS'd584409367, `RNS_PRIME_BITS'd128504548, `RNS_PRIME_BITS'd1198110666, `RNS_PRIME_BITS'd2093525380, `RNS_PRIME_BITS'd1018779229},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd2069863598, `RNS_PRIME_BITS'd393295591, `RNS_PRIME_BITS'd662574108, `RNS_PRIME_BITS'd1618984568, `RNS_PRIME_BITS'd1897061504, `RNS_PRIME_BITS'd1626894753, `RNS_PRIME_BITS'd785660546, `RNS_PRIME_BITS'd1741429703, `RNS_PRIME_BITS'd1351549263, `RNS_PRIME_BITS'd175983492},
			'{`RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd213582633, `RNS_PRIME_BITS'd357115202, `RNS_PRIME_BITS'd131829033, `RNS_PRIME_BITS'd1912147431, `RNS_PRIME_BITS'd1125024231, `RNS_PRIME_BITS'd112369863, `RNS_PRIME_BITS'd1887587115, `RNS_PRIME_BITS'd172071841, `RNS_PRIME_BITS'd3267222, `RNS_PRIME_BITS'd392999815},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1533865378, `RNS_PRIME_BITS'd1582349081, `RNS_PRIME_BITS'd55207768, `RNS_PRIME_BITS'd982311399, `RNS_PRIME_BITS'd2042751230, `RNS_PRIME_BITS'd1591140899, `RNS_PRIME_BITS'd1977620904, `RNS_PRIME_BITS'd1151693408, `RNS_PRIME_BITS'd962289971, `RNS_PRIME_BITS'd1216299653},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd1088633814, `RNS_PRIME_BITS'd1620652108, `RNS_PRIME_BITS'd1072859780, `RNS_PRIME_BITS'd1716492589, `RNS_PRIME_BITS'd1878641723, `RNS_PRIME_BITS'd424479118, `RNS_PRIME_BITS'd676148982, `RNS_PRIME_BITS'd1291675146, `RNS_PRIME_BITS'd275045412, `RNS_PRIME_BITS'd2137120005},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1100413384, `RNS_PRIME_BITS'd1978143492, `RNS_PRIME_BITS'd150820397, `RNS_PRIME_BITS'd122126806, `RNS_PRIME_BITS'd805125457, `RNS_PRIME_BITS'd1957598273, `RNS_PRIME_BITS'd1664211415, `RNS_PRIME_BITS'd433820530, `RNS_PRIME_BITS'd1031212423, `RNS_PRIME_BITS'd2075850888},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd455645603, `RNS_PRIME_BITS'd1437973548, `RNS_PRIME_BITS'd526094255, `RNS_PRIME_BITS'd1471406618, `RNS_PRIME_BITS'd626364197, `RNS_PRIME_BITS'd1097850551, `RNS_PRIME_BITS'd283569171, `RNS_PRIME_BITS'd1967627634, `RNS_PRIME_BITS'd629099459, `RNS_PRIME_BITS'd220754807},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd404173944, `RNS_PRIME_BITS'd1280370870, `RNS_PRIME_BITS'd1680036814, `RNS_PRIME_BITS'd831415558, `RNS_PRIME_BITS'd1453466998, `RNS_PRIME_BITS'd1251323311, `RNS_PRIME_BITS'd178595888, `RNS_PRIME_BITS'd1301726056, `RNS_PRIME_BITS'd682894469, `RNS_PRIME_BITS'd998942748},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd1802592268, `RNS_PRIME_BITS'd538562524, `RNS_PRIME_BITS'd754433925, `RNS_PRIME_BITS'd758098834, `RNS_PRIME_BITS'd508378035, `RNS_PRIME_BITS'd16158829, `RNS_PRIME_BITS'd398410764, `RNS_PRIME_BITS'd1323421910, `RNS_PRIME_BITS'd574860302, `RNS_PRIME_BITS'd230198794},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1298870339, `RNS_PRIME_BITS'd1371966331, `RNS_PRIME_BITS'd486775603, `RNS_PRIME_BITS'd1745595608, `RNS_PRIME_BITS'd977139072, `RNS_PRIME_BITS'd1577615387, `RNS_PRIME_BITS'd845388841, `RNS_PRIME_BITS'd1383409292, `RNS_PRIME_BITS'd1156098269, `RNS_PRIME_BITS'd511049232},
			'{`RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd776469658, `RNS_PRIME_BITS'd868886789, `RNS_PRIME_BITS'd1111228649, `RNS_PRIME_BITS'd1682930164, `RNS_PRIME_BITS'd1482616654, `RNS_PRIME_BITS'd19795401, `RNS_PRIME_BITS'd916066367, `RNS_PRIME_BITS'd410369712, `RNS_PRIME_BITS'd1508628942, `RNS_PRIME_BITS'd1027616005},
			'{`RNS_PRIME_BITS'd65, `RNS_PRIME_BITS'd288608023, `RNS_PRIME_BITS'd884875679, `RNS_PRIME_BITS'd2129793745, `RNS_PRIME_BITS'd1390612102, `RNS_PRIME_BITS'd1247469495, `RNS_PRIME_BITS'd402421964, `RNS_PRIME_BITS'd171389492, `RNS_PRIME_BITS'd847018695, `RNS_PRIME_BITS'd423659366, `RNS_PRIME_BITS'd306751802},
			'{`RNS_PRIME_BITS'd125, `RNS_PRIME_BITS'd1400454688, `RNS_PRIME_BITS'd458343670, `RNS_PRIME_BITS'd1676856052, `RNS_PRIME_BITS'd1547931005, `RNS_PRIME_BITS'd1672360936, `RNS_PRIME_BITS'd1294908542, `RNS_PRIME_BITS'd1883743919, `RNS_PRIME_BITS'd1902095418, `RNS_PRIME_BITS'd863501120, `RNS_PRIME_BITS'd1528679881},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd1432061567, `RNS_PRIME_BITS'd1049079374, `RNS_PRIME_BITS'd1799349082, `RNS_PRIME_BITS'd79483802, `RNS_PRIME_BITS'd1345695708, `RNS_PRIME_BITS'd906954780, `RNS_PRIME_BITS'd270142736, `RNS_PRIME_BITS'd192165409, `RNS_PRIME_BITS'd875758123, `RNS_PRIME_BITS'd2086154122},
			'{`RNS_PRIME_BITS'd126, `RNS_PRIME_BITS'd403126479, `RNS_PRIME_BITS'd560593487, `RNS_PRIME_BITS'd2130249107, `RNS_PRIME_BITS'd685480156, `RNS_PRIME_BITS'd531025128, `RNS_PRIME_BITS'd1961020752, `RNS_PRIME_BITS'd1416004345, `RNS_PRIME_BITS'd1163312518, `RNS_PRIME_BITS'd542940595, `RNS_PRIME_BITS'd1602361313},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd1876170776, `RNS_PRIME_BITS'd207817282, `RNS_PRIME_BITS'd1845188263, `RNS_PRIME_BITS'd718249832, `RNS_PRIME_BITS'd1560307015, `RNS_PRIME_BITS'd2062247605, `RNS_PRIME_BITS'd1295592290, `RNS_PRIME_BITS'd182989956, `RNS_PRIME_BITS'd1039082331, `RNS_PRIME_BITS'd1004878744},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1322405792, `RNS_PRIME_BITS'd447313531, `RNS_PRIME_BITS'd1237321093, `RNS_PRIME_BITS'd1836164500, `RNS_PRIME_BITS'd967516334, `RNS_PRIME_BITS'd1969034683, `RNS_PRIME_BITS'd224303424, `RNS_PRIME_BITS'd1204719006, `RNS_PRIME_BITS'd501510025, `RNS_PRIME_BITS'd449478465},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1800622512, `RNS_PRIME_BITS'd11502919, `RNS_PRIME_BITS'd1359284997, `RNS_PRIME_BITS'd1554821509, `RNS_PRIME_BITS'd1368860510, `RNS_PRIME_BITS'd1515534217, `RNS_PRIME_BITS'd853345787, `RNS_PRIME_BITS'd898890556, `RNS_PRIME_BITS'd438314314, `RNS_PRIME_BITS'd314609344},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd539995158, `RNS_PRIME_BITS'd1100988721, `RNS_PRIME_BITS'd1569959951, `RNS_PRIME_BITS'd487920310, `RNS_PRIME_BITS'd1006328958, `RNS_PRIME_BITS'd162787508, `RNS_PRIME_BITS'd1814019566, `RNS_PRIME_BITS'd832497277, `RNS_PRIME_BITS'd599188777, `RNS_PRIME_BITS'd937650948},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd1338848872, `RNS_PRIME_BITS'd605295099, `RNS_PRIME_BITS'd452374042, `RNS_PRIME_BITS'd1445773540, `RNS_PRIME_BITS'd1486283427, `RNS_PRIME_BITS'd2069473118, `RNS_PRIME_BITS'd374373251, `RNS_PRIME_BITS'd1741624734, `RNS_PRIME_BITS'd348229676, `RNS_PRIME_BITS'd1774419076},
			'{`RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd1905201961, `RNS_PRIME_BITS'd1901826682, `RNS_PRIME_BITS'd77363047, `RNS_PRIME_BITS'd1061093330, `RNS_PRIME_BITS'd870546618, `RNS_PRIME_BITS'd39360310, `RNS_PRIME_BITS'd245997636, `RNS_PRIME_BITS'd643896956, `RNS_PRIME_BITS'd589540382, `RNS_PRIME_BITS'd1028180016},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd1520530191, `RNS_PRIME_BITS'd1755924718, `RNS_PRIME_BITS'd914285141, `RNS_PRIME_BITS'd1759093381, `RNS_PRIME_BITS'd234690810, `RNS_PRIME_BITS'd840599770, `RNS_PRIME_BITS'd2026019051, `RNS_PRIME_BITS'd1371268095, `RNS_PRIME_BITS'd1668969470, `RNS_PRIME_BITS'd1575294654},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1350355407, `RNS_PRIME_BITS'd585365704, `RNS_PRIME_BITS'd102464309, `RNS_PRIME_BITS'd161406928, `RNS_PRIME_BITS'd399782264, `RNS_PRIME_BITS'd2092395771, `RNS_PRIME_BITS'd1379603410, `RNS_PRIME_BITS'd43747838, `RNS_PRIME_BITS'd2033233595, `RNS_PRIME_BITS'd787496917},
			'{`RNS_PRIME_BITS'd204, `RNS_PRIME_BITS'd758919575, `RNS_PRIME_BITS'd1038714162, `RNS_PRIME_BITS'd241657437, `RNS_PRIME_BITS'd1656514028, `RNS_PRIME_BITS'd1910945911, `RNS_PRIME_BITS'd1494617399, `RNS_PRIME_BITS'd1212535367, `RNS_PRIME_BITS'd1728632934, `RNS_PRIME_BITS'd985423930, `RNS_PRIME_BITS'd538814506},
			'{`RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd540790257, `RNS_PRIME_BITS'd282549950, `RNS_PRIME_BITS'd1102971969, `RNS_PRIME_BITS'd178205439, `RNS_PRIME_BITS'd204048911, `RNS_PRIME_BITS'd1760218867, `RNS_PRIME_BITS'd218752685, `RNS_PRIME_BITS'd1952199074, `RNS_PRIME_BITS'd528412527, `RNS_PRIME_BITS'd1361892571}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd1200080509, `RNS_PRIME_BITS'd763442823, `RNS_PRIME_BITS'd1484820538, `RNS_PRIME_BITS'd1346537126, `RNS_PRIME_BITS'd474639971, `RNS_PRIME_BITS'd1212249536, `RNS_PRIME_BITS'd1242393698, `RNS_PRIME_BITS'd202839496, `RNS_PRIME_BITS'd1206162087, `RNS_PRIME_BITS'd828332497},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd891524214, `RNS_PRIME_BITS'd1333330448, `RNS_PRIME_BITS'd937730223, `RNS_PRIME_BITS'd1930730694, `RNS_PRIME_BITS'd1647871677, `RNS_PRIME_BITS'd1423732290, `RNS_PRIME_BITS'd188338168, `RNS_PRIME_BITS'd1014250624, `RNS_PRIME_BITS'd151687182, `RNS_PRIME_BITS'd1675291255},
			'{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd822597495, `RNS_PRIME_BITS'd397553203, `RNS_PRIME_BITS'd1195311369, `RNS_PRIME_BITS'd1647793094, `RNS_PRIME_BITS'd1972592422, `RNS_PRIME_BITS'd830420551, `RNS_PRIME_BITS'd1306171775, `RNS_PRIME_BITS'd1717007452, `RNS_PRIME_BITS'd1336192069, `RNS_PRIME_BITS'd728302459},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1570057444, `RNS_PRIME_BITS'd881214540, `RNS_PRIME_BITS'd335677260, `RNS_PRIME_BITS'd1289919525, `RNS_PRIME_BITS'd2004991653, `RNS_PRIME_BITS'd535675211, `RNS_PRIME_BITS'd1350323588, `RNS_PRIME_BITS'd688777921, `RNS_PRIME_BITS'd461933933, `RNS_PRIME_BITS'd1461997536},
			'{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd2081674052, `RNS_PRIME_BITS'd1378730455, `RNS_PRIME_BITS'd1448978258, `RNS_PRIME_BITS'd934481419, `RNS_PRIME_BITS'd1793178076, `RNS_PRIME_BITS'd985866890, `RNS_PRIME_BITS'd1916681940, `RNS_PRIME_BITS'd2119944576, `RNS_PRIME_BITS'd1763992070, `RNS_PRIME_BITS'd1671691132},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd919383396, `RNS_PRIME_BITS'd1469181313, `RNS_PRIME_BITS'd2128218561, `RNS_PRIME_BITS'd1058786009, `RNS_PRIME_BITS'd1617117485, `RNS_PRIME_BITS'd1977676637, `RNS_PRIME_BITS'd760672768, `RNS_PRIME_BITS'd926320549, `RNS_PRIME_BITS'd645779785, `RNS_PRIME_BITS'd1723306563},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd223364879, `RNS_PRIME_BITS'd1101959303, `RNS_PRIME_BITS'd1289088672, `RNS_PRIME_BITS'd28224519, `RNS_PRIME_BITS'd359774853, `RNS_PRIME_BITS'd420855412, `RNS_PRIME_BITS'd1998280500, `RNS_PRIME_BITS'd617091063, `RNS_PRIME_BITS'd1844958825, `RNS_PRIME_BITS'd763414480},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd1236482082, `RNS_PRIME_BITS'd1628826831, `RNS_PRIME_BITS'd2014332492, `RNS_PRIME_BITS'd2145397032, `RNS_PRIME_BITS'd891324508, `RNS_PRIME_BITS'd127235876, `RNS_PRIME_BITS'd650232187, `RNS_PRIME_BITS'd1078749484, `RNS_PRIME_BITS'd1880847675, `RNS_PRIME_BITS'd104270828},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd2105851821, `RNS_PRIME_BITS'd1296491484, `RNS_PRIME_BITS'd640318528, `RNS_PRIME_BITS'd101181268, `RNS_PRIME_BITS'd1804061973, `RNS_PRIME_BITS'd1155373511, `RNS_PRIME_BITS'd403778980, `RNS_PRIME_BITS'd2005259638, `RNS_PRIME_BITS'd1405079551, `RNS_PRIME_BITS'd1043269760},
			'{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd163525889, `RNS_PRIME_BITS'd912265790, `RNS_PRIME_BITS'd1973055876, `RNS_PRIME_BITS'd1498720147, `RNS_PRIME_BITS'd212846886, `RNS_PRIME_BITS'd840146082, `RNS_PRIME_BITS'd400523254, `RNS_PRIME_BITS'd279546007, `RNS_PRIME_BITS'd686680337, `RNS_PRIME_BITS'd921334185},
			'{`RNS_PRIME_BITS'd91, `RNS_PRIME_BITS'd2062015611, `RNS_PRIME_BITS'd49505889, `RNS_PRIME_BITS'd303440329, `RNS_PRIME_BITS'd66022722, `RNS_PRIME_BITS'd563643546, `RNS_PRIME_BITS'd2072257897, `RNS_PRIME_BITS'd2073078718, `RNS_PRIME_BITS'd37105287, `RNS_PRIME_BITS'd1271947553, `RNS_PRIME_BITS'd1977072030},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd970815792, `RNS_PRIME_BITS'd192707806, `RNS_PRIME_BITS'd1141308600, `RNS_PRIME_BITS'd1477484913, `RNS_PRIME_BITS'd43176284, `RNS_PRIME_BITS'd1316492366, `RNS_PRIME_BITS'd1182934014, `RNS_PRIME_BITS'd1662309201, `RNS_PRIME_BITS'd1041752332, `RNS_PRIME_BITS'd1218105870},
			'{`RNS_PRIME_BITS'd230, `RNS_PRIME_BITS'd2003497983, `RNS_PRIME_BITS'd1958520665, `RNS_PRIME_BITS'd371065667, `RNS_PRIME_BITS'd1819481174, `RNS_PRIME_BITS'd1473188219, `RNS_PRIME_BITS'd1037894696, `RNS_PRIME_BITS'd934074797, `RNS_PRIME_BITS'd1239041895, `RNS_PRIME_BITS'd1018626605, `RNS_PRIME_BITS'd1833274154},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd193487518, `RNS_PRIME_BITS'd1513279713, `RNS_PRIME_BITS'd1420062902, `RNS_PRIME_BITS'd827351316, `RNS_PRIME_BITS'd496954541, `RNS_PRIME_BITS'd876760657, `RNS_PRIME_BITS'd382771808, `RNS_PRIME_BITS'd1124157171, `RNS_PRIME_BITS'd260255897, `RNS_PRIME_BITS'd1485252797},
			'{`RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd633840958, `RNS_PRIME_BITS'd607958266, `RNS_PRIME_BITS'd1456860445, `RNS_PRIME_BITS'd1148791822, `RNS_PRIME_BITS'd1899162940, `RNS_PRIME_BITS'd1714832292, `RNS_PRIME_BITS'd164538465, `RNS_PRIME_BITS'd1678588811, `RNS_PRIME_BITS'd1991925171, `RNS_PRIME_BITS'd453252111},
			'{`RNS_PRIME_BITS'd190, `RNS_PRIME_BITS'd467191868, `RNS_PRIME_BITS'd759612476, `RNS_PRIME_BITS'd756111247, `RNS_PRIME_BITS'd1541282745, `RNS_PRIME_BITS'd1206656270, `RNS_PRIME_BITS'd47755363, `RNS_PRIME_BITS'd1444882251, `RNS_PRIME_BITS'd1677771737, `RNS_PRIME_BITS'd848286553, `RNS_PRIME_BITS'd90675889},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd2008979584, `RNS_PRIME_BITS'd1180998593, `RNS_PRIME_BITS'd1057316779, `RNS_PRIME_BITS'd145821606, `RNS_PRIME_BITS'd1360712491, `RNS_PRIME_BITS'd124651113, `RNS_PRIME_BITS'd434741380, `RNS_PRIME_BITS'd192163496, `RNS_PRIME_BITS'd768900022, `RNS_PRIME_BITS'd1526892344},
			'{`RNS_PRIME_BITS'd12, `RNS_PRIME_BITS'd1734286468, `RNS_PRIME_BITS'd1588493249, `RNS_PRIME_BITS'd1298309805, `RNS_PRIME_BITS'd1849929261, `RNS_PRIME_BITS'd750495499, `RNS_PRIME_BITS'd625023951, `RNS_PRIME_BITS'd220893203, `RNS_PRIME_BITS'd1706738073, `RNS_PRIME_BITS'd508176396, `RNS_PRIME_BITS'd4555031},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd948012605, `RNS_PRIME_BITS'd1196284155, `RNS_PRIME_BITS'd550797531, `RNS_PRIME_BITS'd851474140, `RNS_PRIME_BITS'd129815228, `RNS_PRIME_BITS'd866923202, `RNS_PRIME_BITS'd1421302811, `RNS_PRIME_BITS'd1393406885, `RNS_PRIME_BITS'd1666548817, `RNS_PRIME_BITS'd1128831632},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd1774475899, `RNS_PRIME_BITS'd569257811, `RNS_PRIME_BITS'd152504836, `RNS_PRIME_BITS'd2101480885, `RNS_PRIME_BITS'd1641953187, `RNS_PRIME_BITS'd174760499, `RNS_PRIME_BITS'd1548762735, `RNS_PRIME_BITS'd423243704, `RNS_PRIME_BITS'd1645991948, `RNS_PRIME_BITS'd14670732},
			'{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd412839743, `RNS_PRIME_BITS'd2061056607, `RNS_PRIME_BITS'd1665480578, `RNS_PRIME_BITS'd1104325974, `RNS_PRIME_BITS'd1683362402, `RNS_PRIME_BITS'd1840827861, `RNS_PRIME_BITS'd1502220019, `RNS_PRIME_BITS'd958811398, `RNS_PRIME_BITS'd1874827467, `RNS_PRIME_BITS'd739536953},
			'{`RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd1630713082, `RNS_PRIME_BITS'd1263954710, `RNS_PRIME_BITS'd1163208817, `RNS_PRIME_BITS'd1216114114, `RNS_PRIME_BITS'd613916439, `RNS_PRIME_BITS'd1942884202, `RNS_PRIME_BITS'd1456710070, `RNS_PRIME_BITS'd2034850846, `RNS_PRIME_BITS'd1789891369, `RNS_PRIME_BITS'd1164586761},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1025470468, `RNS_PRIME_BITS'd1464807210, `RNS_PRIME_BITS'd26926476, `RNS_PRIME_BITS'd684382674, `RNS_PRIME_BITS'd320027528, `RNS_PRIME_BITS'd175272615, `RNS_PRIME_BITS'd2126398942, `RNS_PRIME_BITS'd1180212133, `RNS_PRIME_BITS'd638731105, `RNS_PRIME_BITS'd1282754145},
			'{`RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd1209988830, `RNS_PRIME_BITS'd1813810395, `RNS_PRIME_BITS'd1443851282, `RNS_PRIME_BITS'd1014522755, `RNS_PRIME_BITS'd1794194528, `RNS_PRIME_BITS'd1499867222, `RNS_PRIME_BITS'd104849238, `RNS_PRIME_BITS'd664868333, `RNS_PRIME_BITS'd844839718, `RNS_PRIME_BITS'd885387120},
			'{`RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd960187279, `RNS_PRIME_BITS'd653992228, `RNS_PRIME_BITS'd1761999657, `RNS_PRIME_BITS'd1926077813, `RNS_PRIME_BITS'd639542810, `RNS_PRIME_BITS'd1118070023, `RNS_PRIME_BITS'd36559994, `RNS_PRIME_BITS'd401381791, `RNS_PRIME_BITS'd1474103760, `RNS_PRIME_BITS'd1154000673},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1516683545, `RNS_PRIME_BITS'd2058751455, `RNS_PRIME_BITS'd1784367478, `RNS_PRIME_BITS'd1851303057, `RNS_PRIME_BITS'd429093524, `RNS_PRIME_BITS'd965831999, `RNS_PRIME_BITS'd921530196, `RNS_PRIME_BITS'd424834983, `RNS_PRIME_BITS'd537392815, `RNS_PRIME_BITS'd1790938327},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd590639415, `RNS_PRIME_BITS'd1116703056, `RNS_PRIME_BITS'd1662792900, `RNS_PRIME_BITS'd325374409, `RNS_PRIME_BITS'd1968431154, `RNS_PRIME_BITS'd938907122, `RNS_PRIME_BITS'd2116561545, `RNS_PRIME_BITS'd1941657490, `RNS_PRIME_BITS'd1415497784, `RNS_PRIME_BITS'd803889223},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd1384648831, `RNS_PRIME_BITS'd1704920161, `RNS_PRIME_BITS'd1473286404, `RNS_PRIME_BITS'd1137006988, `RNS_PRIME_BITS'd646478039, `RNS_PRIME_BITS'd514729890, `RNS_PRIME_BITS'd1407792314, `RNS_PRIME_BITS'd1647232733, `RNS_PRIME_BITS'd487215355, `RNS_PRIME_BITS'd1537506574},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd439141142, `RNS_PRIME_BITS'd1105554982, `RNS_PRIME_BITS'd321560694, `RNS_PRIME_BITS'd1215438488, `RNS_PRIME_BITS'd1135159611, `RNS_PRIME_BITS'd1506584845, `RNS_PRIME_BITS'd647493572, `RNS_PRIME_BITS'd343328089, `RNS_PRIME_BITS'd573750136, `RNS_PRIME_BITS'd800429863},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd1976463683, `RNS_PRIME_BITS'd132410604, `RNS_PRIME_BITS'd1144255464, `RNS_PRIME_BITS'd216961108, `RNS_PRIME_BITS'd267802614, `RNS_PRIME_BITS'd1769983617, `RNS_PRIME_BITS'd1820208699, `RNS_PRIME_BITS'd953884582, `RNS_PRIME_BITS'd429295120, `RNS_PRIME_BITS'd2039157456},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd52698100, `RNS_PRIME_BITS'd1285918303, `RNS_PRIME_BITS'd1357566287, `RNS_PRIME_BITS'd1875655475, `RNS_PRIME_BITS'd1883152018, `RNS_PRIME_BITS'd1280110543, `RNS_PRIME_BITS'd755707142, `RNS_PRIME_BITS'd51240376, `RNS_PRIME_BITS'd784061208, `RNS_PRIME_BITS'd499238714},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd2115348719, `RNS_PRIME_BITS'd1629553037, `RNS_PRIME_BITS'd2090126794, `RNS_PRIME_BITS'd1876890492, `RNS_PRIME_BITS'd1573038377, `RNS_PRIME_BITS'd647548685, `RNS_PRIME_BITS'd1749076506, `RNS_PRIME_BITS'd945220220, `RNS_PRIME_BITS'd1918737536, `RNS_PRIME_BITS'd717973590},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1525932444, `RNS_PRIME_BITS'd673791377, `RNS_PRIME_BITS'd970519012, `RNS_PRIME_BITS'd1654670461, `RNS_PRIME_BITS'd61311357, `RNS_PRIME_BITS'd765335506, `RNS_PRIME_BITS'd1905971639, `RNS_PRIME_BITS'd89398820, `RNS_PRIME_BITS'd461188950, `RNS_PRIME_BITS'd1804005868},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd432244941, `RNS_PRIME_BITS'd1976493473, `RNS_PRIME_BITS'd1420438061, `RNS_PRIME_BITS'd159058146, `RNS_PRIME_BITS'd93482918, `RNS_PRIME_BITS'd1529264452, `RNS_PRIME_BITS'd1224842106, `RNS_PRIME_BITS'd1799131946, `RNS_PRIME_BITS'd1148288630, `RNS_PRIME_BITS'd1342939113},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd1631643541, `RNS_PRIME_BITS'd172712982, `RNS_PRIME_BITS'd1457337220, `RNS_PRIME_BITS'd1748605590, `RNS_PRIME_BITS'd46778378, `RNS_PRIME_BITS'd470506969, `RNS_PRIME_BITS'd2137214118, `RNS_PRIME_BITS'd1157468964, `RNS_PRIME_BITS'd1360670059, `RNS_PRIME_BITS'd229065900},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1618976126, `RNS_PRIME_BITS'd1904130676, `RNS_PRIME_BITS'd1819072910, `RNS_PRIME_BITS'd1756297114, `RNS_PRIME_BITS'd1866884845, `RNS_PRIME_BITS'd26246128, `RNS_PRIME_BITS'd1456488456, `RNS_PRIME_BITS'd1161703571, `RNS_PRIME_BITS'd715811823, `RNS_PRIME_BITS'd116577021},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd1899595082, `RNS_PRIME_BITS'd1278318011, `RNS_PRIME_BITS'd271800990, `RNS_PRIME_BITS'd1514842438, `RNS_PRIME_BITS'd1828229785, `RNS_PRIME_BITS'd2113377357, `RNS_PRIME_BITS'd194612482, `RNS_PRIME_BITS'd156633970, `RNS_PRIME_BITS'd1423913066, `RNS_PRIME_BITS'd518914533},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd1844278566, `RNS_PRIME_BITS'd2137593196, `RNS_PRIME_BITS'd973806648, `RNS_PRIME_BITS'd1707162045, `RNS_PRIME_BITS'd1334387408, `RNS_PRIME_BITS'd1308604994, `RNS_PRIME_BITS'd517085582, `RNS_PRIME_BITS'd1407457352, `RNS_PRIME_BITS'd983357796, `RNS_PRIME_BITS'd281358814},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd1937473937, `RNS_PRIME_BITS'd1638713913, `RNS_PRIME_BITS'd1311956334, `RNS_PRIME_BITS'd401395652, `RNS_PRIME_BITS'd1166445832, `RNS_PRIME_BITS'd2105309178, `RNS_PRIME_BITS'd1881755709, `RNS_PRIME_BITS'd1194012134, `RNS_PRIME_BITS'd1491738860, `RNS_PRIME_BITS'd2027617542},
			'{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd211811947, `RNS_PRIME_BITS'd2101772780, `RNS_PRIME_BITS'd777669155, `RNS_PRIME_BITS'd1434645721, `RNS_PRIME_BITS'd583994698, `RNS_PRIME_BITS'd1506977633, `RNS_PRIME_BITS'd348687923, `RNS_PRIME_BITS'd1413294812, `RNS_PRIME_BITS'd1313478566, `RNS_PRIME_BITS'd2050163644},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd962918169, `RNS_PRIME_BITS'd638025505, `RNS_PRIME_BITS'd724515655, `RNS_PRIME_BITS'd1815795451, `RNS_PRIME_BITS'd1238507799, `RNS_PRIME_BITS'd1396565994, `RNS_PRIME_BITS'd1912626561, `RNS_PRIME_BITS'd595609515, `RNS_PRIME_BITS'd1545166810, `RNS_PRIME_BITS'd1569739340},
			'{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd1339421014, `RNS_PRIME_BITS'd30860741, `RNS_PRIME_BITS'd510460971, `RNS_PRIME_BITS'd452478694, `RNS_PRIME_BITS'd1116051042, `RNS_PRIME_BITS'd1200695789, `RNS_PRIME_BITS'd1654999026, `RNS_PRIME_BITS'd2083716470, `RNS_PRIME_BITS'd32485612, `RNS_PRIME_BITS'd2043898978},
			'{`RNS_PRIME_BITS'd65, `RNS_PRIME_BITS'd457488461, `RNS_PRIME_BITS'd957385022, `RNS_PRIME_BITS'd720190009, `RNS_PRIME_BITS'd2112386252, `RNS_PRIME_BITS'd1281451491, `RNS_PRIME_BITS'd255418271, `RNS_PRIME_BITS'd2105666848, `RNS_PRIME_BITS'd2081360100, `RNS_PRIME_BITS'd106491746, `RNS_PRIME_BITS'd573071827},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd458871321, `RNS_PRIME_BITS'd1730557423, `RNS_PRIME_BITS'd556366691, `RNS_PRIME_BITS'd609820826, `RNS_PRIME_BITS'd20629794, `RNS_PRIME_BITS'd621784114, `RNS_PRIME_BITS'd64425472, `RNS_PRIME_BITS'd1318280939, `RNS_PRIME_BITS'd1684336806, `RNS_PRIME_BITS'd342144954},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd1863873852, `RNS_PRIME_BITS'd1872438510, `RNS_PRIME_BITS'd921087366, `RNS_PRIME_BITS'd2144644878, `RNS_PRIME_BITS'd27020329, `RNS_PRIME_BITS'd855233046, `RNS_PRIME_BITS'd851695226, `RNS_PRIME_BITS'd352336188, `RNS_PRIME_BITS'd1416067201, `RNS_PRIME_BITS'd1268747797},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd283443916, `RNS_PRIME_BITS'd1721226539, `RNS_PRIME_BITS'd833625170, `RNS_PRIME_BITS'd2126046509, `RNS_PRIME_BITS'd1899224924, `RNS_PRIME_BITS'd560410923, `RNS_PRIME_BITS'd638363327, `RNS_PRIME_BITS'd979166170, `RNS_PRIME_BITS'd1393182292, `RNS_PRIME_BITS'd998559205},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd1090917356, `RNS_PRIME_BITS'd546170396, `RNS_PRIME_BITS'd541987875, `RNS_PRIME_BITS'd1656918860, `RNS_PRIME_BITS'd1129481157, `RNS_PRIME_BITS'd1558198545, `RNS_PRIME_BITS'd1405374861, `RNS_PRIME_BITS'd630366127, `RNS_PRIME_BITS'd18582012, `RNS_PRIME_BITS'd325595908},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd186953147, `RNS_PRIME_BITS'd1082267987, `RNS_PRIME_BITS'd636419231, `RNS_PRIME_BITS'd453151562, `RNS_PRIME_BITS'd925709971, `RNS_PRIME_BITS'd1970173601, `RNS_PRIME_BITS'd601555226, `RNS_PRIME_BITS'd1372966187, `RNS_PRIME_BITS'd1096191258, `RNS_PRIME_BITS'd1888927148},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd2027719036, `RNS_PRIME_BITS'd1944257985, `RNS_PRIME_BITS'd1488632368, `RNS_PRIME_BITS'd2032677459, `RNS_PRIME_BITS'd1143964994, `RNS_PRIME_BITS'd1778026114, `RNS_PRIME_BITS'd709446183, `RNS_PRIME_BITS'd784025088, `RNS_PRIME_BITS'd1692178668, `RNS_PRIME_BITS'd773383831},
			'{`RNS_PRIME_BITS'd172, `RNS_PRIME_BITS'd439018481, `RNS_PRIME_BITS'd211371316, `RNS_PRIME_BITS'd2039161619, `RNS_PRIME_BITS'd1646244420, `RNS_PRIME_BITS'd1405385353, `RNS_PRIME_BITS'd410277524, `RNS_PRIME_BITS'd219168354, `RNS_PRIME_BITS'd2097150821, `RNS_PRIME_BITS'd249621367, `RNS_PRIME_BITS'd213267524},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd1899645327, `RNS_PRIME_BITS'd1033132759, `RNS_PRIME_BITS'd569691229, `RNS_PRIME_BITS'd2086602616, `RNS_PRIME_BITS'd965989769, `RNS_PRIME_BITS'd1218904279, `RNS_PRIME_BITS'd164520117, `RNS_PRIME_BITS'd841236770, `RNS_PRIME_BITS'd1625608693, `RNS_PRIME_BITS'd2110432411},
			'{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd612885219, `RNS_PRIME_BITS'd871852656, `RNS_PRIME_BITS'd403827737, `RNS_PRIME_BITS'd1680996266, `RNS_PRIME_BITS'd736993401, `RNS_PRIME_BITS'd965118418, `RNS_PRIME_BITS'd479991442, `RNS_PRIME_BITS'd1824998840, `RNS_PRIME_BITS'd5169436, `RNS_PRIME_BITS'd748004077},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd444057103, `RNS_PRIME_BITS'd2131255240, `RNS_PRIME_BITS'd66062368, `RNS_PRIME_BITS'd934030232, `RNS_PRIME_BITS'd242818288, `RNS_PRIME_BITS'd1570700407, `RNS_PRIME_BITS'd541197374, `RNS_PRIME_BITS'd2018139923, `RNS_PRIME_BITS'd1614077085, `RNS_PRIME_BITS'd1593093262},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd1612263438, `RNS_PRIME_BITS'd1971430824, `RNS_PRIME_BITS'd38755249, `RNS_PRIME_BITS'd1995194677, `RNS_PRIME_BITS'd200522088, `RNS_PRIME_BITS'd582810395, `RNS_PRIME_BITS'd1266966648, `RNS_PRIME_BITS'd344688967, `RNS_PRIME_BITS'd1060213806, `RNS_PRIME_BITS'd2023561018},
			'{`RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd1812996810, `RNS_PRIME_BITS'd957282495, `RNS_PRIME_BITS'd121563201, `RNS_PRIME_BITS'd2080312906, `RNS_PRIME_BITS'd1169944814, `RNS_PRIME_BITS'd1685311202, `RNS_PRIME_BITS'd923506844, `RNS_PRIME_BITS'd1393733270, `RNS_PRIME_BITS'd192408217, `RNS_PRIME_BITS'd1399864864},
			'{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd785603745, `RNS_PRIME_BITS'd1124985575, `RNS_PRIME_BITS'd615333184, `RNS_PRIME_BITS'd171239065, `RNS_PRIME_BITS'd917716939, `RNS_PRIME_BITS'd379422610, `RNS_PRIME_BITS'd1131541075, `RNS_PRIME_BITS'd132357192, `RNS_PRIME_BITS'd531028801, `RNS_PRIME_BITS'd2099801308},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd666962800, `RNS_PRIME_BITS'd626395948, `RNS_PRIME_BITS'd2129396256, `RNS_PRIME_BITS'd225107080, `RNS_PRIME_BITS'd1773691326, `RNS_PRIME_BITS'd106636344, `RNS_PRIME_BITS'd1310382114, `RNS_PRIME_BITS'd1357670501, `RNS_PRIME_BITS'd1395505153, `RNS_PRIME_BITS'd1598777259},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd414279160, `RNS_PRIME_BITS'd2105132443, `RNS_PRIME_BITS'd1319820234, `RNS_PRIME_BITS'd1940354682, `RNS_PRIME_BITS'd1671155681, `RNS_PRIME_BITS'd1276229235, `RNS_PRIME_BITS'd1087497670, `RNS_PRIME_BITS'd1366930064, `RNS_PRIME_BITS'd1065288050, `RNS_PRIME_BITS'd789514090},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd676935856, `RNS_PRIME_BITS'd66246684, `RNS_PRIME_BITS'd98329321, `RNS_PRIME_BITS'd758645852, `RNS_PRIME_BITS'd2025924581, `RNS_PRIME_BITS'd1121354722, `RNS_PRIME_BITS'd392540516, `RNS_PRIME_BITS'd1984433100, `RNS_PRIME_BITS'd1374195933, `RNS_PRIME_BITS'd1435123857},
			'{`RNS_PRIME_BITS'd227, `RNS_PRIME_BITS'd371234096, `RNS_PRIME_BITS'd1787218782, `RNS_PRIME_BITS'd1701045119, `RNS_PRIME_BITS'd1315707994, `RNS_PRIME_BITS'd1635389272, `RNS_PRIME_BITS'd1537517337, `RNS_PRIME_BITS'd164586667, `RNS_PRIME_BITS'd767755665, `RNS_PRIME_BITS'd1406324977, `RNS_PRIME_BITS'd421707839},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd794783012, `RNS_PRIME_BITS'd1826476315, `RNS_PRIME_BITS'd745073070, `RNS_PRIME_BITS'd61161766, `RNS_PRIME_BITS'd1626202944, `RNS_PRIME_BITS'd697389653, `RNS_PRIME_BITS'd462336964, `RNS_PRIME_BITS'd613405372, `RNS_PRIME_BITS'd516570002, `RNS_PRIME_BITS'd259736751},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd29260770, `RNS_PRIME_BITS'd1737627983, `RNS_PRIME_BITS'd1368869236, `RNS_PRIME_BITS'd87001412, `RNS_PRIME_BITS'd751321334, `RNS_PRIME_BITS'd1630449349, `RNS_PRIME_BITS'd1925009020, `RNS_PRIME_BITS'd165895353, `RNS_PRIME_BITS'd1757323816, `RNS_PRIME_BITS'd1981692589},
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd1651456045, `RNS_PRIME_BITS'd777036710, `RNS_PRIME_BITS'd913974786, `RNS_PRIME_BITS'd443761781, `RNS_PRIME_BITS'd843980992, `RNS_PRIME_BITS'd108659671, `RNS_PRIME_BITS'd69882638, `RNS_PRIME_BITS'd523247484, `RNS_PRIME_BITS'd859832927, `RNS_PRIME_BITS'd1531594590},
			'{`RNS_PRIME_BITS'd190, `RNS_PRIME_BITS'd107136460, `RNS_PRIME_BITS'd1331473365, `RNS_PRIME_BITS'd1296117632, `RNS_PRIME_BITS'd464633907, `RNS_PRIME_BITS'd1732414836, `RNS_PRIME_BITS'd1578948057, `RNS_PRIME_BITS'd1101251283, `RNS_PRIME_BITS'd953571006, `RNS_PRIME_BITS'd1142589435, `RNS_PRIME_BITS'd941194445}
		},
		'{
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1009470868, `RNS_PRIME_BITS'd1059285696, `RNS_PRIME_BITS'd2111233726, `RNS_PRIME_BITS'd1181797225, `RNS_PRIME_BITS'd247281365, `RNS_PRIME_BITS'd1361098303, `RNS_PRIME_BITS'd123358107, `RNS_PRIME_BITS'd242562007, `RNS_PRIME_BITS'd615074991, `RNS_PRIME_BITS'd863066751},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd1442526389, `RNS_PRIME_BITS'd1451109765, `RNS_PRIME_BITS'd759570929, `RNS_PRIME_BITS'd967366892, `RNS_PRIME_BITS'd1150400084, `RNS_PRIME_BITS'd15337751, `RNS_PRIME_BITS'd1159036390, `RNS_PRIME_BITS'd349349524, `RNS_PRIME_BITS'd1163012136, `RNS_PRIME_BITS'd465414601},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd750152803, `RNS_PRIME_BITS'd1829933038, `RNS_PRIME_BITS'd1493823543, `RNS_PRIME_BITS'd1875110396, `RNS_PRIME_BITS'd1801125890, `RNS_PRIME_BITS'd1439413401, `RNS_PRIME_BITS'd1742873227, `RNS_PRIME_BITS'd670511588, `RNS_PRIME_BITS'd1747943317, `RNS_PRIME_BITS'd1041121805},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd710667216, `RNS_PRIME_BITS'd668291911, `RNS_PRIME_BITS'd1551590314, `RNS_PRIME_BITS'd1336834785, `RNS_PRIME_BITS'd1444222809, `RNS_PRIME_BITS'd1289706156, `RNS_PRIME_BITS'd263459150, `RNS_PRIME_BITS'd787782833, `RNS_PRIME_BITS'd1297067852, `RNS_PRIME_BITS'd763707720},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd462333545, `RNS_PRIME_BITS'd164908801, `RNS_PRIME_BITS'd1359208565, `RNS_PRIME_BITS'd27965648, `RNS_PRIME_BITS'd1300046472, `RNS_PRIME_BITS'd2067187695, `RNS_PRIME_BITS'd2003620841, `RNS_PRIME_BITS'd68295893, `RNS_PRIME_BITS'd393596632, `RNS_PRIME_BITS'd1531113603},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd29321032, `RNS_PRIME_BITS'd182575421, `RNS_PRIME_BITS'd278767608, `RNS_PRIME_BITS'd13039238, `RNS_PRIME_BITS'd125387399, `RNS_PRIME_BITS'd866362783, `RNS_PRIME_BITS'd546754785, `RNS_PRIME_BITS'd1444534331, `RNS_PRIME_BITS'd1890925428, `RNS_PRIME_BITS'd398507953},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd776072300, `RNS_PRIME_BITS'd369934971, `RNS_PRIME_BITS'd227758919, `RNS_PRIME_BITS'd663782441, `RNS_PRIME_BITS'd458406541, `RNS_PRIME_BITS'd365634198, `RNS_PRIME_BITS'd1646649250, `RNS_PRIME_BITS'd522055818, `RNS_PRIME_BITS'd1536596467, `RNS_PRIME_BITS'd731884929},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd584859687, `RNS_PRIME_BITS'd545558731, `RNS_PRIME_BITS'd1016573244, `RNS_PRIME_BITS'd1952727179, `RNS_PRIME_BITS'd253279305, `RNS_PRIME_BITS'd1334123241, `RNS_PRIME_BITS'd1008700734, `RNS_PRIME_BITS'd1406452731, `RNS_PRIME_BITS'd553709607, `RNS_PRIME_BITS'd2067079290},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd1274320930, `RNS_PRIME_BITS'd1051013682, `RNS_PRIME_BITS'd835137478, `RNS_PRIME_BITS'd940287153, `RNS_PRIME_BITS'd953306789, `RNS_PRIME_BITS'd1378780652, `RNS_PRIME_BITS'd462905938, `RNS_PRIME_BITS'd589158728, `RNS_PRIME_BITS'd409679285, `RNS_PRIME_BITS'd322548258},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1052646347, `RNS_PRIME_BITS'd1783112931, `RNS_PRIME_BITS'd579770387, `RNS_PRIME_BITS'd25783435, `RNS_PRIME_BITS'd714395869, `RNS_PRIME_BITS'd926194220, `RNS_PRIME_BITS'd1042065187, `RNS_PRIME_BITS'd1182875176, `RNS_PRIME_BITS'd772639330, `RNS_PRIME_BITS'd2048512099},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd1188558339, `RNS_PRIME_BITS'd25859123, `RNS_PRIME_BITS'd1402308235, `RNS_PRIME_BITS'd1712754601, `RNS_PRIME_BITS'd1923927322, `RNS_PRIME_BITS'd1624727620, `RNS_PRIME_BITS'd498264284, `RNS_PRIME_BITS'd893420920, `RNS_PRIME_BITS'd712555561, `RNS_PRIME_BITS'd1947319725},
			'{`RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd258614282, `RNS_PRIME_BITS'd1928133435, `RNS_PRIME_BITS'd804465547, `RNS_PRIME_BITS'd1156625053, `RNS_PRIME_BITS'd451939450, `RNS_PRIME_BITS'd1065559142, `RNS_PRIME_BITS'd473803265, `RNS_PRIME_BITS'd1342000381, `RNS_PRIME_BITS'd110110599, `RNS_PRIME_BITS'd1888006177},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd1134151760, `RNS_PRIME_BITS'd1025900155, `RNS_PRIME_BITS'd152616605, `RNS_PRIME_BITS'd1084853198, `RNS_PRIME_BITS'd1587489764, `RNS_PRIME_BITS'd393276416, `RNS_PRIME_BITS'd833206810, `RNS_PRIME_BITS'd1512183846, `RNS_PRIME_BITS'd1107732375, `RNS_PRIME_BITS'd202189896},
			'{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd1986256040, `RNS_PRIME_BITS'd64925176, `RNS_PRIME_BITS'd1897807860, `RNS_PRIME_BITS'd1075519612, `RNS_PRIME_BITS'd2124261292, `RNS_PRIME_BITS'd1522680041, `RNS_PRIME_BITS'd875792708, `RNS_PRIME_BITS'd1024182283, `RNS_PRIME_BITS'd736391371, `RNS_PRIME_BITS'd2025394541},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd1102467797, `RNS_PRIME_BITS'd869705189, `RNS_PRIME_BITS'd982880964, `RNS_PRIME_BITS'd1149887003, `RNS_PRIME_BITS'd1489315964, `RNS_PRIME_BITS'd1594313981, `RNS_PRIME_BITS'd1596741645, `RNS_PRIME_BITS'd47209066, `RNS_PRIME_BITS'd65697955, `RNS_PRIME_BITS'd370647466},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd1454706047, `RNS_PRIME_BITS'd1957089326, `RNS_PRIME_BITS'd2055603187, `RNS_PRIME_BITS'd1984132663, `RNS_PRIME_BITS'd1135649691, `RNS_PRIME_BITS'd1662994161, `RNS_PRIME_BITS'd382738037, `RNS_PRIME_BITS'd1021971747, `RNS_PRIME_BITS'd1278410394, `RNS_PRIME_BITS'd848224197},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1960108574, `RNS_PRIME_BITS'd103380166, `RNS_PRIME_BITS'd765355584, `RNS_PRIME_BITS'd1790343184, `RNS_PRIME_BITS'd1180818787, `RNS_PRIME_BITS'd1315372860, `RNS_PRIME_BITS'd2109955717, `RNS_PRIME_BITS'd1532923695, `RNS_PRIME_BITS'd1923098084, `RNS_PRIME_BITS'd1967163199},
			'{`RNS_PRIME_BITS'd224, `RNS_PRIME_BITS'd1026333312, `RNS_PRIME_BITS'd488247527, `RNS_PRIME_BITS'd1408808103, `RNS_PRIME_BITS'd186924908, `RNS_PRIME_BITS'd2102548236, `RNS_PRIME_BITS'd1685512027, `RNS_PRIME_BITS'd1345139168, `RNS_PRIME_BITS'd665775992, `RNS_PRIME_BITS'd293572954, `RNS_PRIME_BITS'd1044202429},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd350046012, `RNS_PRIME_BITS'd692888927, `RNS_PRIME_BITS'd1289240307, `RNS_PRIME_BITS'd1437965560, `RNS_PRIME_BITS'd1626327539, `RNS_PRIME_BITS'd651499330, `RNS_PRIME_BITS'd1932676579, `RNS_PRIME_BITS'd1769051997, `RNS_PRIME_BITS'd1436050154, `RNS_PRIME_BITS'd1422601932},
			'{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd1251135523, `RNS_PRIME_BITS'd1503054959, `RNS_PRIME_BITS'd1591537956, `RNS_PRIME_BITS'd175875939, `RNS_PRIME_BITS'd686042313, `RNS_PRIME_BITS'd789349359, `RNS_PRIME_BITS'd2061586537, `RNS_PRIME_BITS'd1000174230, `RNS_PRIME_BITS'd1967664296, `RNS_PRIME_BITS'd1166387702},
			'{`RNS_PRIME_BITS'd200, `RNS_PRIME_BITS'd830965375, `RNS_PRIME_BITS'd666344643, `RNS_PRIME_BITS'd1138367538, `RNS_PRIME_BITS'd320577083, `RNS_PRIME_BITS'd1108841302, `RNS_PRIME_BITS'd1578237303, `RNS_PRIME_BITS'd1865739296, `RNS_PRIME_BITS'd725731967, `RNS_PRIME_BITS'd1941393888, `RNS_PRIME_BITS'd928846493},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd1109404577, `RNS_PRIME_BITS'd56077653, `RNS_PRIME_BITS'd487662290, `RNS_PRIME_BITS'd1526036730, `RNS_PRIME_BITS'd218540837, `RNS_PRIME_BITS'd8426645, `RNS_PRIME_BITS'd1724894356, `RNS_PRIME_BITS'd119601129, `RNS_PRIME_BITS'd994885796, `RNS_PRIME_BITS'd679393555},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd701444928, `RNS_PRIME_BITS'd1443650031, `RNS_PRIME_BITS'd592589355, `RNS_PRIME_BITS'd1084072119, `RNS_PRIME_BITS'd246542376, `RNS_PRIME_BITS'd379929266, `RNS_PRIME_BITS'd335854879, `RNS_PRIME_BITS'd1786189421, `RNS_PRIME_BITS'd473927344, `RNS_PRIME_BITS'd471571547},
			'{`RNS_PRIME_BITS'd160, `RNS_PRIME_BITS'd799335563, `RNS_PRIME_BITS'd2117568780, `RNS_PRIME_BITS'd1808342590, `RNS_PRIME_BITS'd1703355604, `RNS_PRIME_BITS'd1489793377, `RNS_PRIME_BITS'd1462471817, `RNS_PRIME_BITS'd62641534, `RNS_PRIME_BITS'd1330720306, `RNS_PRIME_BITS'd228950030, `RNS_PRIME_BITS'd1294756401},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd1280218571, `RNS_PRIME_BITS'd276998317, `RNS_PRIME_BITS'd287241555, `RNS_PRIME_BITS'd55231539, `RNS_PRIME_BITS'd1775884151, `RNS_PRIME_BITS'd452586280, `RNS_PRIME_BITS'd240640897, `RNS_PRIME_BITS'd11753761, `RNS_PRIME_BITS'd238629784, `RNS_PRIME_BITS'd702224878},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd490616979, `RNS_PRIME_BITS'd1257988395, `RNS_PRIME_BITS'd1991574628, `RNS_PRIME_BITS'd1985640119, `RNS_PRIME_BITS'd1988620316, `RNS_PRIME_BITS'd1532492693, `RNS_PRIME_BITS'd722930848, `RNS_PRIME_BITS'd713222110, `RNS_PRIME_BITS'd1315700581, `RNS_PRIME_BITS'd1808474522},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd247659990, `RNS_PRIME_BITS'd1758407913, `RNS_PRIME_BITS'd1694139987, `RNS_PRIME_BITS'd1345840427, `RNS_PRIME_BITS'd918392640, `RNS_PRIME_BITS'd981422668, `RNS_PRIME_BITS'd1526005080, `RNS_PRIME_BITS'd1080601395, `RNS_PRIME_BITS'd1650271623, `RNS_PRIME_BITS'd825298036},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd1361957359, `RNS_PRIME_BITS'd2063185659, `RNS_PRIME_BITS'd496129353, `RNS_PRIME_BITS'd378797372, `RNS_PRIME_BITS'd631696779, `RNS_PRIME_BITS'd728602523, `RNS_PRIME_BITS'd812060380, `RNS_PRIME_BITS'd1670949785, `RNS_PRIME_BITS'd764613510, `RNS_PRIME_BITS'd1068795310},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd900600717, `RNS_PRIME_BITS'd730427235, `RNS_PRIME_BITS'd39320506, `RNS_PRIME_BITS'd343493147, `RNS_PRIME_BITS'd1353547960, `RNS_PRIME_BITS'd686545203, `RNS_PRIME_BITS'd696211803, `RNS_PRIME_BITS'd919769245, `RNS_PRIME_BITS'd390224565, `RNS_PRIME_BITS'd644808198},
			'{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd311704809, `RNS_PRIME_BITS'd719625662, `RNS_PRIME_BITS'd1289951375, `RNS_PRIME_BITS'd829841573, `RNS_PRIME_BITS'd1542148888, `RNS_PRIME_BITS'd367970497, `RNS_PRIME_BITS'd1408347597, `RNS_PRIME_BITS'd1716690743, `RNS_PRIME_BITS'd296856234, `RNS_PRIME_BITS'd808350262},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd758837113, `RNS_PRIME_BITS'd1100329447, `RNS_PRIME_BITS'd368852670, `RNS_PRIME_BITS'd1581735370, `RNS_PRIME_BITS'd1083284991, `RNS_PRIME_BITS'd145442452, `RNS_PRIME_BITS'd837745832, `RNS_PRIME_BITS'd484100261, `RNS_PRIME_BITS'd1414331751, `RNS_PRIME_BITS'd2070023642},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd498540477, `RNS_PRIME_BITS'd1866791845, `RNS_PRIME_BITS'd1416227655, `RNS_PRIME_BITS'd1898845419, `RNS_PRIME_BITS'd1310515840, `RNS_PRIME_BITS'd1814212182, `RNS_PRIME_BITS'd622370869, `RNS_PRIME_BITS'd772693883, `RNS_PRIME_BITS'd510090006, `RNS_PRIME_BITS'd1305547028},
			'{`RNS_PRIME_BITS'd140, `RNS_PRIME_BITS'd1546649576, `RNS_PRIME_BITS'd895286725, `RNS_PRIME_BITS'd842210869, `RNS_PRIME_BITS'd1561090691, `RNS_PRIME_BITS'd1834519240, `RNS_PRIME_BITS'd1296221727, `RNS_PRIME_BITS'd1502974055, `RNS_PRIME_BITS'd1279951733, `RNS_PRIME_BITS'd368539140, `RNS_PRIME_BITS'd1928117067},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd1029539639, `RNS_PRIME_BITS'd661360835, `RNS_PRIME_BITS'd878566878, `RNS_PRIME_BITS'd74117403, `RNS_PRIME_BITS'd1932822312, `RNS_PRIME_BITS'd1689401371, `RNS_PRIME_BITS'd1719878186, `RNS_PRIME_BITS'd663073079, `RNS_PRIME_BITS'd17650418, `RNS_PRIME_BITS'd2050149540},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1296344853, `RNS_PRIME_BITS'd597501113, `RNS_PRIME_BITS'd2131263730, `RNS_PRIME_BITS'd1379536769, `RNS_PRIME_BITS'd1025851230, `RNS_PRIME_BITS'd725601243, `RNS_PRIME_BITS'd1686662972, `RNS_PRIME_BITS'd369307577, `RNS_PRIME_BITS'd2111023232, `RNS_PRIME_BITS'd1141517862},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd1437340160, `RNS_PRIME_BITS'd149454194, `RNS_PRIME_BITS'd448800502, `RNS_PRIME_BITS'd634087985, `RNS_PRIME_BITS'd2023115971, `RNS_PRIME_BITS'd47785983, `RNS_PRIME_BITS'd1637028686, `RNS_PRIME_BITS'd1958321872, `RNS_PRIME_BITS'd1089077457, `RNS_PRIME_BITS'd485532887},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd1472077975, `RNS_PRIME_BITS'd1974461403, `RNS_PRIME_BITS'd919247806, `RNS_PRIME_BITS'd122740397, `RNS_PRIME_BITS'd1731404142, `RNS_PRIME_BITS'd1473896036, `RNS_PRIME_BITS'd1199552215, `RNS_PRIME_BITS'd1700085192, `RNS_PRIME_BITS'd2144994216, `RNS_PRIME_BITS'd1448788264},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd529375206, `RNS_PRIME_BITS'd1162201192, `RNS_PRIME_BITS'd1049271176, `RNS_PRIME_BITS'd714619438, `RNS_PRIME_BITS'd507380745, `RNS_PRIME_BITS'd1682110858, `RNS_PRIME_BITS'd149153493, `RNS_PRIME_BITS'd495285705, `RNS_PRIME_BITS'd195140134, `RNS_PRIME_BITS'd7931349},
			'{`RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd1747753193, `RNS_PRIME_BITS'd808639625, `RNS_PRIME_BITS'd472538066, `RNS_PRIME_BITS'd1571339800, `RNS_PRIME_BITS'd1654261788, `RNS_PRIME_BITS'd705175539, `RNS_PRIME_BITS'd1708906822, `RNS_PRIME_BITS'd2001809947, `RNS_PRIME_BITS'd1566405094, `RNS_PRIME_BITS'd2100156635},
			'{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd1552215765, `RNS_PRIME_BITS'd1517289410, `RNS_PRIME_BITS'd740138996, `RNS_PRIME_BITS'd1330230427, `RNS_PRIME_BITS'd800086174, `RNS_PRIME_BITS'd853088201, `RNS_PRIME_BITS'd1751615510, `RNS_PRIME_BITS'd816071205, `RNS_PRIME_BITS'd457182357, `RNS_PRIME_BITS'd117971729},
			'{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd334073626, `RNS_PRIME_BITS'd325426827, `RNS_PRIME_BITS'd338529955, `RNS_PRIME_BITS'd1266845221, `RNS_PRIME_BITS'd2135109857, `RNS_PRIME_BITS'd1663552532, `RNS_PRIME_BITS'd1248351113, `RNS_PRIME_BITS'd1290182204, `RNS_PRIME_BITS'd1477367240, `RNS_PRIME_BITS'd124667059},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1830954722, `RNS_PRIME_BITS'd77711468, `RNS_PRIME_BITS'd700385416, `RNS_PRIME_BITS'd948951932, `RNS_PRIME_BITS'd2028309788, `RNS_PRIME_BITS'd1240393211, `RNS_PRIME_BITS'd951719519, `RNS_PRIME_BITS'd135667951, `RNS_PRIME_BITS'd547064396, `RNS_PRIME_BITS'd380839980},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd745827786, `RNS_PRIME_BITS'd1298707808, `RNS_PRIME_BITS'd1600423691, `RNS_PRIME_BITS'd1666779003, `RNS_PRIME_BITS'd220829526, `RNS_PRIME_BITS'd1240770819, `RNS_PRIME_BITS'd1685187343, `RNS_PRIME_BITS'd2120946560, `RNS_PRIME_BITS'd710020422, `RNS_PRIME_BITS'd815915178},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd617001839, `RNS_PRIME_BITS'd721997401, `RNS_PRIME_BITS'd1518924378, `RNS_PRIME_BITS'd1590096494, `RNS_PRIME_BITS'd1842965493, `RNS_PRIME_BITS'd147797285, `RNS_PRIME_BITS'd99377221, `RNS_PRIME_BITS'd1940338333, `RNS_PRIME_BITS'd1183061368, `RNS_PRIME_BITS'd55939493},
			'{`RNS_PRIME_BITS'd109, `RNS_PRIME_BITS'd1781673816, `RNS_PRIME_BITS'd1660080103, `RNS_PRIME_BITS'd675151357, `RNS_PRIME_BITS'd284839445, `RNS_PRIME_BITS'd1721630828, `RNS_PRIME_BITS'd929351696, `RNS_PRIME_BITS'd648747942, `RNS_PRIME_BITS'd1441319413, `RNS_PRIME_BITS'd147403764, `RNS_PRIME_BITS'd894500788},
			'{`RNS_PRIME_BITS'd167, `RNS_PRIME_BITS'd1638764536, `RNS_PRIME_BITS'd226155562, `RNS_PRIME_BITS'd1558965399, `RNS_PRIME_BITS'd1652348663, `RNS_PRIME_BITS'd183477659, `RNS_PRIME_BITS'd1240445966, `RNS_PRIME_BITS'd1378172289, `RNS_PRIME_BITS'd964968083, `RNS_PRIME_BITS'd1434266727, `RNS_PRIME_BITS'd1949960722},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd892621167, `RNS_PRIME_BITS'd715403974, `RNS_PRIME_BITS'd1667342200, `RNS_PRIME_BITS'd1850572720, `RNS_PRIME_BITS'd1448992807, `RNS_PRIME_BITS'd693728774, `RNS_PRIME_BITS'd1436366742, `RNS_PRIME_BITS'd218246604, `RNS_PRIME_BITS'd99657321, `RNS_PRIME_BITS'd1484284312},
			'{`RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd471980412, `RNS_PRIME_BITS'd85841037, `RNS_PRIME_BITS'd1806989352, `RNS_PRIME_BITS'd839662003, `RNS_PRIME_BITS'd204365264, `RNS_PRIME_BITS'd902788342, `RNS_PRIME_BITS'd1629482838, `RNS_PRIME_BITS'd761710908, `RNS_PRIME_BITS'd1553042948, `RNS_PRIME_BITS'd1370346074},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd395248194, `RNS_PRIME_BITS'd508633201, `RNS_PRIME_BITS'd1003648148, `RNS_PRIME_BITS'd742960557, `RNS_PRIME_BITS'd1199934404, `RNS_PRIME_BITS'd1140683490, `RNS_PRIME_BITS'd2070623744, `RNS_PRIME_BITS'd1009812673, `RNS_PRIME_BITS'd1517003674, `RNS_PRIME_BITS'd1854109449},
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd197675820, `RNS_PRIME_BITS'd1553414174, `RNS_PRIME_BITS'd1363601577, `RNS_PRIME_BITS'd877727289, `RNS_PRIME_BITS'd778884704, `RNS_PRIME_BITS'd140765190, `RNS_PRIME_BITS'd824461665, `RNS_PRIME_BITS'd338628839, `RNS_PRIME_BITS'd1864591341, `RNS_PRIME_BITS'd1034729952},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd639052355, `RNS_PRIME_BITS'd1724638488, `RNS_PRIME_BITS'd256578571, `RNS_PRIME_BITS'd2042373287, `RNS_PRIME_BITS'd1976228615, `RNS_PRIME_BITS'd1329985515, `RNS_PRIME_BITS'd608129761, `RNS_PRIME_BITS'd1062540116, `RNS_PRIME_BITS'd827546522, `RNS_PRIME_BITS'd643207208},
			'{`RNS_PRIME_BITS'd38, `RNS_PRIME_BITS'd173839089, `RNS_PRIME_BITS'd623443047, `RNS_PRIME_BITS'd2081485343, `RNS_PRIME_BITS'd2021888097, `RNS_PRIME_BITS'd1895098558, `RNS_PRIME_BITS'd1356856977, `RNS_PRIME_BITS'd196006464, `RNS_PRIME_BITS'd1515332419, `RNS_PRIME_BITS'd1417149033, `RNS_PRIME_BITS'd649886345},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd1599165080, `RNS_PRIME_BITS'd1519620434, `RNS_PRIME_BITS'd991407211, `RNS_PRIME_BITS'd1683409177, `RNS_PRIME_BITS'd218342411, `RNS_PRIME_BITS'd1221308268, `RNS_PRIME_BITS'd505773069, `RNS_PRIME_BITS'd508555322, `RNS_PRIME_BITS'd2136420968, `RNS_PRIME_BITS'd810470118},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd215500260, `RNS_PRIME_BITS'd708429966, `RNS_PRIME_BITS'd1001171908, `RNS_PRIME_BITS'd1072297728, `RNS_PRIME_BITS'd585730913, `RNS_PRIME_BITS'd406587165, `RNS_PRIME_BITS'd1403067124, `RNS_PRIME_BITS'd71420301, `RNS_PRIME_BITS'd740313291, `RNS_PRIME_BITS'd67466789},
			'{`RNS_PRIME_BITS'd126, `RNS_PRIME_BITS'd828238587, `RNS_PRIME_BITS'd1928339913, `RNS_PRIME_BITS'd1861171605, `RNS_PRIME_BITS'd448561050, `RNS_PRIME_BITS'd775409091, `RNS_PRIME_BITS'd782098569, `RNS_PRIME_BITS'd1156880857, `RNS_PRIME_BITS'd690479185, `RNS_PRIME_BITS'd90001041, `RNS_PRIME_BITS'd1931543640},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd489085046, `RNS_PRIME_BITS'd1733645683, `RNS_PRIME_BITS'd156429143, `RNS_PRIME_BITS'd632607053, `RNS_PRIME_BITS'd1657040578, `RNS_PRIME_BITS'd1173112666, `RNS_PRIME_BITS'd722953706, `RNS_PRIME_BITS'd896254897, `RNS_PRIME_BITS'd918693399, `RNS_PRIME_BITS'd51188377},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd1733374276, `RNS_PRIME_BITS'd2056079262, `RNS_PRIME_BITS'd685988363, `RNS_PRIME_BITS'd2092783309, `RNS_PRIME_BITS'd1124326565, `RNS_PRIME_BITS'd130517758, `RNS_PRIME_BITS'd683747068, `RNS_PRIME_BITS'd1017686349, `RNS_PRIME_BITS'd101652713, `RNS_PRIME_BITS'd968057452},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd907706794, `RNS_PRIME_BITS'd1486913609, `RNS_PRIME_BITS'd169771980, `RNS_PRIME_BITS'd1000920908, `RNS_PRIME_BITS'd1292267408, `RNS_PRIME_BITS'd1503566491, `RNS_PRIME_BITS'd1298860174, `RNS_PRIME_BITS'd1403996731, `RNS_PRIME_BITS'd1495193766, `RNS_PRIME_BITS'd1792685184},
			'{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd142790292, `RNS_PRIME_BITS'd1501961768, `RNS_PRIME_BITS'd1096113647, `RNS_PRIME_BITS'd59008586, `RNS_PRIME_BITS'd547126228, `RNS_PRIME_BITS'd578161108, `RNS_PRIME_BITS'd1342013353, `RNS_PRIME_BITS'd1642049005, `RNS_PRIME_BITS'd1255356727, `RNS_PRIME_BITS'd2022814391},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd1561935038, `RNS_PRIME_BITS'd2017906891, `RNS_PRIME_BITS'd1351345065, `RNS_PRIME_BITS'd381633742, `RNS_PRIME_BITS'd365293597, `RNS_PRIME_BITS'd1402165682, `RNS_PRIME_BITS'd1146911705, `RNS_PRIME_BITS'd366987110, `RNS_PRIME_BITS'd1488630248, `RNS_PRIME_BITS'd235128430},
			'{`RNS_PRIME_BITS'd209, `RNS_PRIME_BITS'd1084494995, `RNS_PRIME_BITS'd1545708908, `RNS_PRIME_BITS'd30256148, `RNS_PRIME_BITS'd451912908, `RNS_PRIME_BITS'd313097157, `RNS_PRIME_BITS'd686155994, `RNS_PRIME_BITS'd556580487, `RNS_PRIME_BITS'd1999485434, `RNS_PRIME_BITS'd1076694426, `RNS_PRIME_BITS'd129794887},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd898750319, `RNS_PRIME_BITS'd172964496, `RNS_PRIME_BITS'd1087776049, `RNS_PRIME_BITS'd1913349342, `RNS_PRIME_BITS'd1119245976, `RNS_PRIME_BITS'd719523378, `RNS_PRIME_BITS'd388986068, `RNS_PRIME_BITS'd184644838, `RNS_PRIME_BITS'd897332067, `RNS_PRIME_BITS'd1477574188},
			'{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd1051762018, `RNS_PRIME_BITS'd963471866, `RNS_PRIME_BITS'd1395442869, `RNS_PRIME_BITS'd358623576, `RNS_PRIME_BITS'd948053553, `RNS_PRIME_BITS'd1005908302, `RNS_PRIME_BITS'd117102706, `RNS_PRIME_BITS'd2127796116, `RNS_PRIME_BITS'd251021151, `RNS_PRIME_BITS'd1689035947},
			'{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd1638282365, `RNS_PRIME_BITS'd2078370330, `RNS_PRIME_BITS'd2071528343, `RNS_PRIME_BITS'd288829682, `RNS_PRIME_BITS'd781078892, `RNS_PRIME_BITS'd1346577202, `RNS_PRIME_BITS'd1254628064, `RNS_PRIME_BITS'd2102459133, `RNS_PRIME_BITS'd1190998108, `RNS_PRIME_BITS'd1056433499}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd98, `RNS_PRIME_BITS'd756944296, `RNS_PRIME_BITS'd122705213, `RNS_PRIME_BITS'd215098579, `RNS_PRIME_BITS'd558880560, `RNS_PRIME_BITS'd1539899998, `RNS_PRIME_BITS'd289848963, `RNS_PRIME_BITS'd1678538925, `RNS_PRIME_BITS'd394191171, `RNS_PRIME_BITS'd634069679, `RNS_PRIME_BITS'd808546167},
			'{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd920288642, `RNS_PRIME_BITS'd619929400, `RNS_PRIME_BITS'd2102004370, `RNS_PRIME_BITS'd658060701, `RNS_PRIME_BITS'd801396733, `RNS_PRIME_BITS'd912877126, `RNS_PRIME_BITS'd590802778, `RNS_PRIME_BITS'd1612507353, `RNS_PRIME_BITS'd864197842, `RNS_PRIME_BITS'd1001485960},
			'{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd348561088, `RNS_PRIME_BITS'd491076128, `RNS_PRIME_BITS'd714422051, `RNS_PRIME_BITS'd1824980246, `RNS_PRIME_BITS'd1284201570, `RNS_PRIME_BITS'd639402279, `RNS_PRIME_BITS'd934641060, `RNS_PRIME_BITS'd403112053, `RNS_PRIME_BITS'd441430335, `RNS_PRIME_BITS'd374077436},
			'{`RNS_PRIME_BITS'd224, `RNS_PRIME_BITS'd1481129075, `RNS_PRIME_BITS'd1173261677, `RNS_PRIME_BITS'd542584225, `RNS_PRIME_BITS'd826233829, `RNS_PRIME_BITS'd424755671, `RNS_PRIME_BITS'd1976301337, `RNS_PRIME_BITS'd1703871749, `RNS_PRIME_BITS'd2058966166, `RNS_PRIME_BITS'd1045314142, `RNS_PRIME_BITS'd444784763},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd2078157161, `RNS_PRIME_BITS'd1086464892, `RNS_PRIME_BITS'd75875424, `RNS_PRIME_BITS'd498481576, `RNS_PRIME_BITS'd1731763468, `RNS_PRIME_BITS'd281387541, `RNS_PRIME_BITS'd219216850, `RNS_PRIME_BITS'd1181602597, `RNS_PRIME_BITS'd332024981, `RNS_PRIME_BITS'd1970123655},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd766104215, `RNS_PRIME_BITS'd897761974, `RNS_PRIME_BITS'd956076791, `RNS_PRIME_BITS'd103025663, `RNS_PRIME_BITS'd413598930, `RNS_PRIME_BITS'd1777119412, `RNS_PRIME_BITS'd62010798, `RNS_PRIME_BITS'd871648428, `RNS_PRIME_BITS'd243525864, `RNS_PRIME_BITS'd53729226},
			'{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd892576806, `RNS_PRIME_BITS'd363204569, `RNS_PRIME_BITS'd146552122, `RNS_PRIME_BITS'd966409010, `RNS_PRIME_BITS'd1181458793, `RNS_PRIME_BITS'd77955920, `RNS_PRIME_BITS'd301653627, `RNS_PRIME_BITS'd887007953, `RNS_PRIME_BITS'd2046375383, `RNS_PRIME_BITS'd2031701742},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1923261626, `RNS_PRIME_BITS'd1626643301, `RNS_PRIME_BITS'd514979862, `RNS_PRIME_BITS'd1692696516, `RNS_PRIME_BITS'd1542994472, `RNS_PRIME_BITS'd1095179054, `RNS_PRIME_BITS'd1479276592, `RNS_PRIME_BITS'd870335140, `RNS_PRIME_BITS'd1447744458, `RNS_PRIME_BITS'd1610026542},
			'{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd1496934724, `RNS_PRIME_BITS'd1799027417, `RNS_PRIME_BITS'd772125838, `RNS_PRIME_BITS'd623108326, `RNS_PRIME_BITS'd162544118, `RNS_PRIME_BITS'd1044467904, `RNS_PRIME_BITS'd123165166, `RNS_PRIME_BITS'd112301653, `RNS_PRIME_BITS'd1885796526, `RNS_PRIME_BITS'd47304881},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1292384931, `RNS_PRIME_BITS'd1283125350, `RNS_PRIME_BITS'd946685954, `RNS_PRIME_BITS'd1566774911, `RNS_PRIME_BITS'd289366889, `RNS_PRIME_BITS'd562482578, `RNS_PRIME_BITS'd755678131, `RNS_PRIME_BITS'd939575002, `RNS_PRIME_BITS'd406787976, `RNS_PRIME_BITS'd1648253748},
			'{`RNS_PRIME_BITS'd250, `RNS_PRIME_BITS'd2041909279, `RNS_PRIME_BITS'd1010644888, `RNS_PRIME_BITS'd237640070, `RNS_PRIME_BITS'd1760368693, `RNS_PRIME_BITS'd1589740421, `RNS_PRIME_BITS'd926878210, `RNS_PRIME_BITS'd333360489, `RNS_PRIME_BITS'd1165931589, `RNS_PRIME_BITS'd381600443, `RNS_PRIME_BITS'd726734272},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1517079098, `RNS_PRIME_BITS'd1644382541, `RNS_PRIME_BITS'd1027549878, `RNS_PRIME_BITS'd1475581490, `RNS_PRIME_BITS'd1373593971, `RNS_PRIME_BITS'd371840760, `RNS_PRIME_BITS'd1175505197, `RNS_PRIME_BITS'd562869800, `RNS_PRIME_BITS'd132614066, `RNS_PRIME_BITS'd723953081},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1751755894, `RNS_PRIME_BITS'd708522738, `RNS_PRIME_BITS'd2080123633, `RNS_PRIME_BITS'd1193926756, `RNS_PRIME_BITS'd586837643, `RNS_PRIME_BITS'd2069125115, `RNS_PRIME_BITS'd185771928, `RNS_PRIME_BITS'd735448522, `RNS_PRIME_BITS'd2105362418, `RNS_PRIME_BITS'd1682303634},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd977179992, `RNS_PRIME_BITS'd1597614454, `RNS_PRIME_BITS'd330755552, `RNS_PRIME_BITS'd1482174494, `RNS_PRIME_BITS'd58627688, `RNS_PRIME_BITS'd1786982976, `RNS_PRIME_BITS'd1093906567, `RNS_PRIME_BITS'd9821198, `RNS_PRIME_BITS'd1014529391, `RNS_PRIME_BITS'd444959520},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1039177960, `RNS_PRIME_BITS'd759707900, `RNS_PRIME_BITS'd1664949726, `RNS_PRIME_BITS'd1910759276, `RNS_PRIME_BITS'd1506167042, `RNS_PRIME_BITS'd342143880, `RNS_PRIME_BITS'd642648445, `RNS_PRIME_BITS'd438351890, `RNS_PRIME_BITS'd1393434614, `RNS_PRIME_BITS'd1609935322},
			'{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd1091024095, `RNS_PRIME_BITS'd1495309039, `RNS_PRIME_BITS'd1495546415, `RNS_PRIME_BITS'd366854486, `RNS_PRIME_BITS'd1946947073, `RNS_PRIME_BITS'd212257074, `RNS_PRIME_BITS'd727108647, `RNS_PRIME_BITS'd1583102579, `RNS_PRIME_BITS'd940288927, `RNS_PRIME_BITS'd1090179883},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd1180437362, `RNS_PRIME_BITS'd1612106737, `RNS_PRIME_BITS'd1579661372, `RNS_PRIME_BITS'd1066963514, `RNS_PRIME_BITS'd1448771346, `RNS_PRIME_BITS'd1634914117, `RNS_PRIME_BITS'd1463381297, `RNS_PRIME_BITS'd788422671, `RNS_PRIME_BITS'd1356471761, `RNS_PRIME_BITS'd856207391},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd2011692313, `RNS_PRIME_BITS'd2083810482, `RNS_PRIME_BITS'd1011138887, `RNS_PRIME_BITS'd1687773689, `RNS_PRIME_BITS'd2042289377, `RNS_PRIME_BITS'd2136052518, `RNS_PRIME_BITS'd365051888, `RNS_PRIME_BITS'd203763502, `RNS_PRIME_BITS'd689785390, `RNS_PRIME_BITS'd388920039},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd2111959884, `RNS_PRIME_BITS'd637192946, `RNS_PRIME_BITS'd1459777859, `RNS_PRIME_BITS'd2082380365, `RNS_PRIME_BITS'd663522106, `RNS_PRIME_BITS'd1312381297, `RNS_PRIME_BITS'd1468520081, `RNS_PRIME_BITS'd15664384, `RNS_PRIME_BITS'd241185211, `RNS_PRIME_BITS'd900842370},
			'{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd1141321336, `RNS_PRIME_BITS'd623216989, `RNS_PRIME_BITS'd1850831334, `RNS_PRIME_BITS'd632862970, `RNS_PRIME_BITS'd1198103764, `RNS_PRIME_BITS'd350286938, `RNS_PRIME_BITS'd367761564, `RNS_PRIME_BITS'd750453388, `RNS_PRIME_BITS'd948501950, `RNS_PRIME_BITS'd207714458},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd178885166, `RNS_PRIME_BITS'd939373248, `RNS_PRIME_BITS'd1047396252, `RNS_PRIME_BITS'd1418532753, `RNS_PRIME_BITS'd590402488, `RNS_PRIME_BITS'd26388965, `RNS_PRIME_BITS'd1315309724, `RNS_PRIME_BITS'd1940759916, `RNS_PRIME_BITS'd317451626, `RNS_PRIME_BITS'd830556876},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd1190772203, `RNS_PRIME_BITS'd157281526, `RNS_PRIME_BITS'd1064716869, `RNS_PRIME_BITS'd651983791, `RNS_PRIME_BITS'd1946561351, `RNS_PRIME_BITS'd922612769, `RNS_PRIME_BITS'd1427588392, `RNS_PRIME_BITS'd1602395720, `RNS_PRIME_BITS'd179629519, `RNS_PRIME_BITS'd1949172089},
			'{`RNS_PRIME_BITS'd14, `RNS_PRIME_BITS'd1626774197, `RNS_PRIME_BITS'd51112652, `RNS_PRIME_BITS'd1414587661, `RNS_PRIME_BITS'd733302685, `RNS_PRIME_BITS'd1863534766, `RNS_PRIME_BITS'd365980552, `RNS_PRIME_BITS'd1406802060, `RNS_PRIME_BITS'd2125255447, `RNS_PRIME_BITS'd1375466702, `RNS_PRIME_BITS'd752600877},
			'{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd634399691, `RNS_PRIME_BITS'd439731941, `RNS_PRIME_BITS'd139938089, `RNS_PRIME_BITS'd1635101342, `RNS_PRIME_BITS'd534522836, `RNS_PRIME_BITS'd193272054, `RNS_PRIME_BITS'd149409975, `RNS_PRIME_BITS'd109253682, `RNS_PRIME_BITS'd536741572, `RNS_PRIME_BITS'd503812547},
			'{`RNS_PRIME_BITS'd14, `RNS_PRIME_BITS'd1521734925, `RNS_PRIME_BITS'd1995547893, `RNS_PRIME_BITS'd2023622907, `RNS_PRIME_BITS'd2055871111, `RNS_PRIME_BITS'd1208401802, `RNS_PRIME_BITS'd1524250380, `RNS_PRIME_BITS'd914433489, `RNS_PRIME_BITS'd1191326138, `RNS_PRIME_BITS'd1552533845, `RNS_PRIME_BITS'd302104206},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd1649189898, `RNS_PRIME_BITS'd1860664494, `RNS_PRIME_BITS'd1587681563, `RNS_PRIME_BITS'd1442017150, `RNS_PRIME_BITS'd924940724, `RNS_PRIME_BITS'd766251788, `RNS_PRIME_BITS'd1366986849, `RNS_PRIME_BITS'd832945064, `RNS_PRIME_BITS'd1438883388, `RNS_PRIME_BITS'd2048972688},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd1430439926, `RNS_PRIME_BITS'd711864433, `RNS_PRIME_BITS'd424322243, `RNS_PRIME_BITS'd418923343, `RNS_PRIME_BITS'd1057817811, `RNS_PRIME_BITS'd872647143, `RNS_PRIME_BITS'd973562595, `RNS_PRIME_BITS'd2079675567, `RNS_PRIME_BITS'd269522458, `RNS_PRIME_BITS'd1158313209},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd1483324892, `RNS_PRIME_BITS'd828872810, `RNS_PRIME_BITS'd634503179, `RNS_PRIME_BITS'd1902772888, `RNS_PRIME_BITS'd1345345209, `RNS_PRIME_BITS'd270898593, `RNS_PRIME_BITS'd393197840, `RNS_PRIME_BITS'd1306138847, `RNS_PRIME_BITS'd800560867, `RNS_PRIME_BITS'd566755435},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd1035863888, `RNS_PRIME_BITS'd169302177, `RNS_PRIME_BITS'd1051655177, `RNS_PRIME_BITS'd72029532, `RNS_PRIME_BITS'd578051517, `RNS_PRIME_BITS'd2020064322, `RNS_PRIME_BITS'd769615588, `RNS_PRIME_BITS'd1415775, `RNS_PRIME_BITS'd1026375119, `RNS_PRIME_BITS'd1624416478},
			'{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd1068378451, `RNS_PRIME_BITS'd2142634691, `RNS_PRIME_BITS'd2023385312, `RNS_PRIME_BITS'd1629040001, `RNS_PRIME_BITS'd288612142, `RNS_PRIME_BITS'd48392507, `RNS_PRIME_BITS'd2031474988, `RNS_PRIME_BITS'd968533341, `RNS_PRIME_BITS'd1708314575, `RNS_PRIME_BITS'd1603721881},
			'{`RNS_PRIME_BITS'd19, `RNS_PRIME_BITS'd1805901599, `RNS_PRIME_BITS'd635588413, `RNS_PRIME_BITS'd674619357, `RNS_PRIME_BITS'd1928671780, `RNS_PRIME_BITS'd1313529070, `RNS_PRIME_BITS'd758454042, `RNS_PRIME_BITS'd1389121571, `RNS_PRIME_BITS'd449356471, `RNS_PRIME_BITS'd1393990720, `RNS_PRIME_BITS'd1411656699},
			'{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd1179149705, `RNS_PRIME_BITS'd651678062, `RNS_PRIME_BITS'd802462086, `RNS_PRIME_BITS'd1433895202, `RNS_PRIME_BITS'd1101101166, `RNS_PRIME_BITS'd1420785745, `RNS_PRIME_BITS'd1453332306, `RNS_PRIME_BITS'd473232344, `RNS_PRIME_BITS'd346011562, `RNS_PRIME_BITS'd362336411},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd128734713, `RNS_PRIME_BITS'd45971329, `RNS_PRIME_BITS'd450357003, `RNS_PRIME_BITS'd430327931, `RNS_PRIME_BITS'd1901081832, `RNS_PRIME_BITS'd1850446329, `RNS_PRIME_BITS'd1356277916, `RNS_PRIME_BITS'd1894009834, `RNS_PRIME_BITS'd1654424258, `RNS_PRIME_BITS'd1389852984},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd1555549702, `RNS_PRIME_BITS'd640145001, `RNS_PRIME_BITS'd55528391, `RNS_PRIME_BITS'd1531193394, `RNS_PRIME_BITS'd1999318179, `RNS_PRIME_BITS'd1980387041, `RNS_PRIME_BITS'd1455622713, `RNS_PRIME_BITS'd337649656, `RNS_PRIME_BITS'd1944971335, `RNS_PRIME_BITS'd39193040},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd615901594, `RNS_PRIME_BITS'd1315420046, `RNS_PRIME_BITS'd661625167, `RNS_PRIME_BITS'd884702839, `RNS_PRIME_BITS'd1092496894, `RNS_PRIME_BITS'd620607668, `RNS_PRIME_BITS'd1158129907, `RNS_PRIME_BITS'd722590365, `RNS_PRIME_BITS'd1743319449, `RNS_PRIME_BITS'd1597766519},
			'{`RNS_PRIME_BITS'd91, `RNS_PRIME_BITS'd450877701, `RNS_PRIME_BITS'd1355462767, `RNS_PRIME_BITS'd1649544237, `RNS_PRIME_BITS'd22741787, `RNS_PRIME_BITS'd1396797963, `RNS_PRIME_BITS'd1513785613, `RNS_PRIME_BITS'd169716184, `RNS_PRIME_BITS'd993672038, `RNS_PRIME_BITS'd997528099, `RNS_PRIME_BITS'd1356980939},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd636514584, `RNS_PRIME_BITS'd106840857, `RNS_PRIME_BITS'd1816193754, `RNS_PRIME_BITS'd872532405, `RNS_PRIME_BITS'd289066761, `RNS_PRIME_BITS'd1162309021, `RNS_PRIME_BITS'd501662822, `RNS_PRIME_BITS'd1275836370, `RNS_PRIME_BITS'd1113616513, `RNS_PRIME_BITS'd1937952304},
			'{`RNS_PRIME_BITS'd227, `RNS_PRIME_BITS'd1349091715, `RNS_PRIME_BITS'd710508274, `RNS_PRIME_BITS'd53916049, `RNS_PRIME_BITS'd892352118, `RNS_PRIME_BITS'd1676317144, `RNS_PRIME_BITS'd68501289, `RNS_PRIME_BITS'd1582074502, `RNS_PRIME_BITS'd990710243, `RNS_PRIME_BITS'd548120542, `RNS_PRIME_BITS'd1503758101},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd1464058483, `RNS_PRIME_BITS'd1876515819, `RNS_PRIME_BITS'd1705897221, `RNS_PRIME_BITS'd630243582, `RNS_PRIME_BITS'd1048021765, `RNS_PRIME_BITS'd2016333840, `RNS_PRIME_BITS'd1214658334, `RNS_PRIME_BITS'd1212061726, `RNS_PRIME_BITS'd435162823, `RNS_PRIME_BITS'd1773298773},
			'{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd672760953, `RNS_PRIME_BITS'd453761589, `RNS_PRIME_BITS'd906525044, `RNS_PRIME_BITS'd1338587845, `RNS_PRIME_BITS'd293737774, `RNS_PRIME_BITS'd1104233153, `RNS_PRIME_BITS'd728564592, `RNS_PRIME_BITS'd1757669185, `RNS_PRIME_BITS'd836311922, `RNS_PRIME_BITS'd1597949330},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd958815012, `RNS_PRIME_BITS'd712388732, `RNS_PRIME_BITS'd1090323550, `RNS_PRIME_BITS'd1401979207, `RNS_PRIME_BITS'd691658176, `RNS_PRIME_BITS'd897853246, `RNS_PRIME_BITS'd130324108, `RNS_PRIME_BITS'd235082293, `RNS_PRIME_BITS'd272908608, `RNS_PRIME_BITS'd1780157505},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd521945284, `RNS_PRIME_BITS'd339461574, `RNS_PRIME_BITS'd426201171, `RNS_PRIME_BITS'd463808127, `RNS_PRIME_BITS'd1117668383, `RNS_PRIME_BITS'd1817644501, `RNS_PRIME_BITS'd269432543, `RNS_PRIME_BITS'd1681520616, `RNS_PRIME_BITS'd1671140741, `RNS_PRIME_BITS'd778800941},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1196318120, `RNS_PRIME_BITS'd943800735, `RNS_PRIME_BITS'd708634853, `RNS_PRIME_BITS'd1275238634, `RNS_PRIME_BITS'd223514494, `RNS_PRIME_BITS'd1301305234, `RNS_PRIME_BITS'd1778337041, `RNS_PRIME_BITS'd1565756285, `RNS_PRIME_BITS'd1567480715, `RNS_PRIME_BITS'd297157374},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1506297267, `RNS_PRIME_BITS'd1044533827, `RNS_PRIME_BITS'd834705683, `RNS_PRIME_BITS'd171373320, `RNS_PRIME_BITS'd1409962622, `RNS_PRIME_BITS'd1084471199, `RNS_PRIME_BITS'd649501518, `RNS_PRIME_BITS'd632785945, `RNS_PRIME_BITS'd238265256, `RNS_PRIME_BITS'd60492361},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd423290649, `RNS_PRIME_BITS'd130161356, `RNS_PRIME_BITS'd433008803, `RNS_PRIME_BITS'd1496588630, `RNS_PRIME_BITS'd205996650, `RNS_PRIME_BITS'd2109215868, `RNS_PRIME_BITS'd1870663145, `RNS_PRIME_BITS'd997244014, `RNS_PRIME_BITS'd820815684, `RNS_PRIME_BITS'd1890365950},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd489118368, `RNS_PRIME_BITS'd53243278, `RNS_PRIME_BITS'd960283879, `RNS_PRIME_BITS'd1370574008, `RNS_PRIME_BITS'd656330380, `RNS_PRIME_BITS'd1213488008, `RNS_PRIME_BITS'd1171567110, `RNS_PRIME_BITS'd2011371095, `RNS_PRIME_BITS'd1450866668, `RNS_PRIME_BITS'd1643834382},
			'{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd1468745573, `RNS_PRIME_BITS'd1500226919, `RNS_PRIME_BITS'd709225644, `RNS_PRIME_BITS'd208641226, `RNS_PRIME_BITS'd1814377724, `RNS_PRIME_BITS'd917546372, `RNS_PRIME_BITS'd247341781, `RNS_PRIME_BITS'd304148312, `RNS_PRIME_BITS'd2005803122, `RNS_PRIME_BITS'd175782463},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd891797542, `RNS_PRIME_BITS'd653086194, `RNS_PRIME_BITS'd768837840, `RNS_PRIME_BITS'd1571602351, `RNS_PRIME_BITS'd2002965606, `RNS_PRIME_BITS'd618366569, `RNS_PRIME_BITS'd767214608, `RNS_PRIME_BITS'd347891498, `RNS_PRIME_BITS'd1840585159, `RNS_PRIME_BITS'd1219775717},
			'{`RNS_PRIME_BITS'd54, `RNS_PRIME_BITS'd1554944681, `RNS_PRIME_BITS'd1945559989, `RNS_PRIME_BITS'd1379795373, `RNS_PRIME_BITS'd779777648, `RNS_PRIME_BITS'd1598838617, `RNS_PRIME_BITS'd1629158868, `RNS_PRIME_BITS'd1173793448, `RNS_PRIME_BITS'd294674157, `RNS_PRIME_BITS'd720406012, `RNS_PRIME_BITS'd1566691276},
			'{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd622292279, `RNS_PRIME_BITS'd894086195, `RNS_PRIME_BITS'd504615667, `RNS_PRIME_BITS'd1267184785, `RNS_PRIME_BITS'd1540570442, `RNS_PRIME_BITS'd2087148003, `RNS_PRIME_BITS'd216383661, `RNS_PRIME_BITS'd2011514501, `RNS_PRIME_BITS'd1832367809, `RNS_PRIME_BITS'd306236817},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1617539343, `RNS_PRIME_BITS'd1509078504, `RNS_PRIME_BITS'd1677255642, `RNS_PRIME_BITS'd1870009396, `RNS_PRIME_BITS'd1219710610, `RNS_PRIME_BITS'd606307754, `RNS_PRIME_BITS'd1776819890, `RNS_PRIME_BITS'd319524168, `RNS_PRIME_BITS'd1374207680, `RNS_PRIME_BITS'd130294610},
			'{`RNS_PRIME_BITS'd188, `RNS_PRIME_BITS'd1067837075, `RNS_PRIME_BITS'd1385439140, `RNS_PRIME_BITS'd659448305, `RNS_PRIME_BITS'd4094954, `RNS_PRIME_BITS'd1089720733, `RNS_PRIME_BITS'd171495281, `RNS_PRIME_BITS'd733383705, `RNS_PRIME_BITS'd1636589514, `RNS_PRIME_BITS'd364098126, `RNS_PRIME_BITS'd387322545},
			'{`RNS_PRIME_BITS'd76, `RNS_PRIME_BITS'd239592500, `RNS_PRIME_BITS'd1254603375, `RNS_PRIME_BITS'd2032032937, `RNS_PRIME_BITS'd429734372, `RNS_PRIME_BITS'd368644292, `RNS_PRIME_BITS'd380403049, `RNS_PRIME_BITS'd353763790, `RNS_PRIME_BITS'd425832415, `RNS_PRIME_BITS'd454966972, `RNS_PRIME_BITS'd858364937},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd621736395, `RNS_PRIME_BITS'd1743918343, `RNS_PRIME_BITS'd953258127, `RNS_PRIME_BITS'd1455230777, `RNS_PRIME_BITS'd1904778140, `RNS_PRIME_BITS'd1725027859, `RNS_PRIME_BITS'd1887240521, `RNS_PRIME_BITS'd953071279, `RNS_PRIME_BITS'd52253894, `RNS_PRIME_BITS'd1396954880},
			'{`RNS_PRIME_BITS'd110, `RNS_PRIME_BITS'd409532192, `RNS_PRIME_BITS'd574621093, `RNS_PRIME_BITS'd1549030169, `RNS_PRIME_BITS'd398031170, `RNS_PRIME_BITS'd1183794060, `RNS_PRIME_BITS'd837754652, `RNS_PRIME_BITS'd357528744, `RNS_PRIME_BITS'd1283685681, `RNS_PRIME_BITS'd147527223, `RNS_PRIME_BITS'd21644912},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd1456289267, `RNS_PRIME_BITS'd1402691139, `RNS_PRIME_BITS'd937558522, `RNS_PRIME_BITS'd980627082, `RNS_PRIME_BITS'd504146054, `RNS_PRIME_BITS'd1197577875, `RNS_PRIME_BITS'd1526814416, `RNS_PRIME_BITS'd1913152867, `RNS_PRIME_BITS'd590089731, `RNS_PRIME_BITS'd313337357},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd715727657, `RNS_PRIME_BITS'd800470511, `RNS_PRIME_BITS'd789514753, `RNS_PRIME_BITS'd29630604, `RNS_PRIME_BITS'd673118526, `RNS_PRIME_BITS'd1964977658, `RNS_PRIME_BITS'd1218860682, `RNS_PRIME_BITS'd443319792, `RNS_PRIME_BITS'd69989357, `RNS_PRIME_BITS'd1171646330},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd803493360, `RNS_PRIME_BITS'd1738387913, `RNS_PRIME_BITS'd304988204, `RNS_PRIME_BITS'd103949306, `RNS_PRIME_BITS'd1502080929, `RNS_PRIME_BITS'd1259467122, `RNS_PRIME_BITS'd1513146771, `RNS_PRIME_BITS'd1710269234, `RNS_PRIME_BITS'd1780488706, `RNS_PRIME_BITS'd2017006981},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd777518755, `RNS_PRIME_BITS'd580980566, `RNS_PRIME_BITS'd1199065696, `RNS_PRIME_BITS'd940006881, `RNS_PRIME_BITS'd2118307795, `RNS_PRIME_BITS'd1943589673, `RNS_PRIME_BITS'd48625062, `RNS_PRIME_BITS'd1847797323, `RNS_PRIME_BITS'd913696679, `RNS_PRIME_BITS'd1313187657},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd888244773, `RNS_PRIME_BITS'd2010020377, `RNS_PRIME_BITS'd1822259321, `RNS_PRIME_BITS'd1363296168, `RNS_PRIME_BITS'd422908440, `RNS_PRIME_BITS'd422263949, `RNS_PRIME_BITS'd421382940, `RNS_PRIME_BITS'd1259006780, `RNS_PRIME_BITS'd2034051697, `RNS_PRIME_BITS'd132281593},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1422934754, `RNS_PRIME_BITS'd320629642, `RNS_PRIME_BITS'd1804652899, `RNS_PRIME_BITS'd560158418, `RNS_PRIME_BITS'd170261745, `RNS_PRIME_BITS'd238064376, `RNS_PRIME_BITS'd567214289, `RNS_PRIME_BITS'd818492995, `RNS_PRIME_BITS'd822408733, `RNS_PRIME_BITS'd189099628},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd170999966, `RNS_PRIME_BITS'd596990475, `RNS_PRIME_BITS'd1124372369, `RNS_PRIME_BITS'd1381310896, `RNS_PRIME_BITS'd1283652987, `RNS_PRIME_BITS'd1815539681, `RNS_PRIME_BITS'd1494873663, `RNS_PRIME_BITS'd1504413265, `RNS_PRIME_BITS'd1509351377, `RNS_PRIME_BITS'd1243923972},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd1079828041, `RNS_PRIME_BITS'd1532609068, `RNS_PRIME_BITS'd2146948539, `RNS_PRIME_BITS'd2059393512, `RNS_PRIME_BITS'd1990753042, `RNS_PRIME_BITS'd1647700813, `RNS_PRIME_BITS'd1570478159, `RNS_PRIME_BITS'd740806793, `RNS_PRIME_BITS'd1397374360, `RNS_PRIME_BITS'd792571087},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd1851629553, `RNS_PRIME_BITS'd817033625, `RNS_PRIME_BITS'd925064124, `RNS_PRIME_BITS'd864472788, `RNS_PRIME_BITS'd2097206050, `RNS_PRIME_BITS'd1180496284, `RNS_PRIME_BITS'd1102888390, `RNS_PRIME_BITS'd1126395253, `RNS_PRIME_BITS'd1730014532, `RNS_PRIME_BITS'd522498877}
		},
		'{
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd2093229614, `RNS_PRIME_BITS'd1594939326, `RNS_PRIME_BITS'd2129408746, `RNS_PRIME_BITS'd515961875, `RNS_PRIME_BITS'd408086754, `RNS_PRIME_BITS'd732875402, `RNS_PRIME_BITS'd2026027002, `RNS_PRIME_BITS'd805570684, `RNS_PRIME_BITS'd1073824354, `RNS_PRIME_BITS'd1510829748},
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd549927883, `RNS_PRIME_BITS'd1670672579, `RNS_PRIME_BITS'd1976836782, `RNS_PRIME_BITS'd210278674, `RNS_PRIME_BITS'd1052894574, `RNS_PRIME_BITS'd567246061, `RNS_PRIME_BITS'd290782795, `RNS_PRIME_BITS'd31825726, `RNS_PRIME_BITS'd22301553, `RNS_PRIME_BITS'd520263245},
			'{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd2052563433, `RNS_PRIME_BITS'd865357411, `RNS_PRIME_BITS'd877206945, `RNS_PRIME_BITS'd332219361, `RNS_PRIME_BITS'd1888000618, `RNS_PRIME_BITS'd492912011, `RNS_PRIME_BITS'd165990016, `RNS_PRIME_BITS'd813220825, `RNS_PRIME_BITS'd773730978, `RNS_PRIME_BITS'd535313993},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd679871904, `RNS_PRIME_BITS'd1391983487, `RNS_PRIME_BITS'd1581918323, `RNS_PRIME_BITS'd6614776, `RNS_PRIME_BITS'd537843598, `RNS_PRIME_BITS'd344276080, `RNS_PRIME_BITS'd215274171, `RNS_PRIME_BITS'd139614015, `RNS_PRIME_BITS'd756993395, `RNS_PRIME_BITS'd1263029922},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd1935986842, `RNS_PRIME_BITS'd297991975, `RNS_PRIME_BITS'd2024739446, `RNS_PRIME_BITS'd1875499490, `RNS_PRIME_BITS'd960656405, `RNS_PRIME_BITS'd1297571181, `RNS_PRIME_BITS'd566473629, `RNS_PRIME_BITS'd1390188342, `RNS_PRIME_BITS'd1167410950, `RNS_PRIME_BITS'd1744004413},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1911044284, `RNS_PRIME_BITS'd1363737647, `RNS_PRIME_BITS'd141726558, `RNS_PRIME_BITS'd1417379962, `RNS_PRIME_BITS'd114365590, `RNS_PRIME_BITS'd1699274536, `RNS_PRIME_BITS'd1923624147, `RNS_PRIME_BITS'd528907992, `RNS_PRIME_BITS'd1358619977, `RNS_PRIME_BITS'd677391043},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd1056493092, `RNS_PRIME_BITS'd979379828, `RNS_PRIME_BITS'd629136779, `RNS_PRIME_BITS'd2042362216, `RNS_PRIME_BITS'd882333075, `RNS_PRIME_BITS'd1645177601, `RNS_PRIME_BITS'd976620806, `RNS_PRIME_BITS'd883773391, `RNS_PRIME_BITS'd217561163, `RNS_PRIME_BITS'd655628344},
			'{`RNS_PRIME_BITS'd172, `RNS_PRIME_BITS'd1302656556, `RNS_PRIME_BITS'd2003565913, `RNS_PRIME_BITS'd2123456021, `RNS_PRIME_BITS'd1319181517, `RNS_PRIME_BITS'd935013258, `RNS_PRIME_BITS'd1315985568, `RNS_PRIME_BITS'd300986754, `RNS_PRIME_BITS'd716833974, `RNS_PRIME_BITS'd1120810093, `RNS_PRIME_BITS'd1359891328},
			'{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd1857983504, `RNS_PRIME_BITS'd740569677, `RNS_PRIME_BITS'd184660302, `RNS_PRIME_BITS'd1437762581, `RNS_PRIME_BITS'd902723789, `RNS_PRIME_BITS'd2032467114, `RNS_PRIME_BITS'd1599659035, `RNS_PRIME_BITS'd1070337855, `RNS_PRIME_BITS'd1250148397, `RNS_PRIME_BITS'd1519553625},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd1895785533, `RNS_PRIME_BITS'd350537742, `RNS_PRIME_BITS'd1889487476, `RNS_PRIME_BITS'd1950941450, `RNS_PRIME_BITS'd1445414645, `RNS_PRIME_BITS'd1203617370, `RNS_PRIME_BITS'd320773000, `RNS_PRIME_BITS'd1640089997, `RNS_PRIME_BITS'd990480866, `RNS_PRIME_BITS'd1307488448},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd189407134, `RNS_PRIME_BITS'd1596578544, `RNS_PRIME_BITS'd1079171263, `RNS_PRIME_BITS'd177257884, `RNS_PRIME_BITS'd1517332314, `RNS_PRIME_BITS'd1856127707, `RNS_PRIME_BITS'd496678922, `RNS_PRIME_BITS'd1471620793, `RNS_PRIME_BITS'd1073270781, `RNS_PRIME_BITS'd54477085},
			'{`RNS_PRIME_BITS'd227, `RNS_PRIME_BITS'd1963677029, `RNS_PRIME_BITS'd1302579369, `RNS_PRIME_BITS'd1949192641, `RNS_PRIME_BITS'd1976665287, `RNS_PRIME_BITS'd1920450121, `RNS_PRIME_BITS'd464648234, `RNS_PRIME_BITS'd291202116, `RNS_PRIME_BITS'd511583183, `RNS_PRIME_BITS'd1574589756, `RNS_PRIME_BITS'd36085905},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd772843475, `RNS_PRIME_BITS'd1251599548, `RNS_PRIME_BITS'd720603763, `RNS_PRIME_BITS'd1115201455, `RNS_PRIME_BITS'd895216401, `RNS_PRIME_BITS'd1759371126, `RNS_PRIME_BITS'd73858778, `RNS_PRIME_BITS'd2101650466, `RNS_PRIME_BITS'd1194696050, `RNS_PRIME_BITS'd1057318020},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd143831775, `RNS_PRIME_BITS'd1335751836, `RNS_PRIME_BITS'd77124490, `RNS_PRIME_BITS'd1724992222, `RNS_PRIME_BITS'd1135294237, `RNS_PRIME_BITS'd1467076272, `RNS_PRIME_BITS'd781303287, `RNS_PRIME_BITS'd703350164, `RNS_PRIME_BITS'd1476954131, `RNS_PRIME_BITS'd1577508282},
			'{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd1563623061, `RNS_PRIME_BITS'd1287843437, `RNS_PRIME_BITS'd2078116520, `RNS_PRIME_BITS'd34615367, `RNS_PRIME_BITS'd403488064, `RNS_PRIME_BITS'd522236936, `RNS_PRIME_BITS'd203328565, `RNS_PRIME_BITS'd2055531390, `RNS_PRIME_BITS'd1662731930, `RNS_PRIME_BITS'd444861306},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd961097731, `RNS_PRIME_BITS'd15364555, `RNS_PRIME_BITS'd1521391975, `RNS_PRIME_BITS'd1802958694, `RNS_PRIME_BITS'd1017961424, `RNS_PRIME_BITS'd1275447412, `RNS_PRIME_BITS'd1469041292, `RNS_PRIME_BITS'd784283701, `RNS_PRIME_BITS'd2129592055, `RNS_PRIME_BITS'd971694289},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd2106140549, `RNS_PRIME_BITS'd466451599, `RNS_PRIME_BITS'd1931916114, `RNS_PRIME_BITS'd1962924317, `RNS_PRIME_BITS'd2047598362, `RNS_PRIME_BITS'd1666192024, `RNS_PRIME_BITS'd1263310145, `RNS_PRIME_BITS'd1650966868, `RNS_PRIME_BITS'd697536728, `RNS_PRIME_BITS'd1521290773},
			'{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd154434647, `RNS_PRIME_BITS'd424742579, `RNS_PRIME_BITS'd1096084947, `RNS_PRIME_BITS'd585866407, `RNS_PRIME_BITS'd2045421985, `RNS_PRIME_BITS'd1366476480, `RNS_PRIME_BITS'd753575197, `RNS_PRIME_BITS'd1106401081, `RNS_PRIME_BITS'd198085369, `RNS_PRIME_BITS'd1348282246},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd1477880774, `RNS_PRIME_BITS'd951624174, `RNS_PRIME_BITS'd760942751, `RNS_PRIME_BITS'd1333811954, `RNS_PRIME_BITS'd136189195, `RNS_PRIME_BITS'd804687059, `RNS_PRIME_BITS'd70250105, `RNS_PRIME_BITS'd1088118474, `RNS_PRIME_BITS'd44726510, `RNS_PRIME_BITS'd172822629},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd528915016, `RNS_PRIME_BITS'd858174682, `RNS_PRIME_BITS'd477590989, `RNS_PRIME_BITS'd1500705855, `RNS_PRIME_BITS'd907451082, `RNS_PRIME_BITS'd998232963, `RNS_PRIME_BITS'd1436084028, `RNS_PRIME_BITS'd2070982410, `RNS_PRIME_BITS'd2125839465, `RNS_PRIME_BITS'd31768294},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd1405848859, `RNS_PRIME_BITS'd1327933209, `RNS_PRIME_BITS'd1841854068, `RNS_PRIME_BITS'd828745487, `RNS_PRIME_BITS'd663100266, `RNS_PRIME_BITS'd1009121487, `RNS_PRIME_BITS'd841510940, `RNS_PRIME_BITS'd52968677, `RNS_PRIME_BITS'd195707468, `RNS_PRIME_BITS'd559310491},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd200746244, `RNS_PRIME_BITS'd162540014, `RNS_PRIME_BITS'd399216368, `RNS_PRIME_BITS'd1691797585, `RNS_PRIME_BITS'd1350310670, `RNS_PRIME_BITS'd1639585619, `RNS_PRIME_BITS'd14514979, `RNS_PRIME_BITS'd1400205831, `RNS_PRIME_BITS'd2054665046, `RNS_PRIME_BITS'd2058034179},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd4796394, `RNS_PRIME_BITS'd2130966831, `RNS_PRIME_BITS'd2013725783, `RNS_PRIME_BITS'd518294556, `RNS_PRIME_BITS'd718697348, `RNS_PRIME_BITS'd1322185413, `RNS_PRIME_BITS'd1808108333, `RNS_PRIME_BITS'd338692487, `RNS_PRIME_BITS'd117530401, `RNS_PRIME_BITS'd1288730022},
			'{`RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd585575613, `RNS_PRIME_BITS'd1554508098, `RNS_PRIME_BITS'd652916945, `RNS_PRIME_BITS'd1058539056, `RNS_PRIME_BITS'd1958584842, `RNS_PRIME_BITS'd1422636540, `RNS_PRIME_BITS'd1100340582, `RNS_PRIME_BITS'd1323900548, `RNS_PRIME_BITS'd1569816373, `RNS_PRIME_BITS'd788198908},
			'{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd344939095, `RNS_PRIME_BITS'd1345453983, `RNS_PRIME_BITS'd2141154022, `RNS_PRIME_BITS'd765958731, `RNS_PRIME_BITS'd1233119841, `RNS_PRIME_BITS'd571343950, `RNS_PRIME_BITS'd740741567, `RNS_PRIME_BITS'd1204512715, `RNS_PRIME_BITS'd1397939535, `RNS_PRIME_BITS'd165909394},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd999767081, `RNS_PRIME_BITS'd113543233, `RNS_PRIME_BITS'd1180636072, `RNS_PRIME_BITS'd525743590, `RNS_PRIME_BITS'd1275760925, `RNS_PRIME_BITS'd2033912442, `RNS_PRIME_BITS'd653197917, `RNS_PRIME_BITS'd6032009, `RNS_PRIME_BITS'd538748257, `RNS_PRIME_BITS'd2021403154},
			'{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd1206089721, `RNS_PRIME_BITS'd175540582, `RNS_PRIME_BITS'd1666691843, `RNS_PRIME_BITS'd96112261, `RNS_PRIME_BITS'd91062146, `RNS_PRIME_BITS'd1619906008, `RNS_PRIME_BITS'd942468398, `RNS_PRIME_BITS'd928366200, `RNS_PRIME_BITS'd1930156748, `RNS_PRIME_BITS'd802807704},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1402637614, `RNS_PRIME_BITS'd1635769260, `RNS_PRIME_BITS'd1060525205, `RNS_PRIME_BITS'd173076347, `RNS_PRIME_BITS'd919279684, `RNS_PRIME_BITS'd863934943, `RNS_PRIME_BITS'd1423614860, `RNS_PRIME_BITS'd1156671880, `RNS_PRIME_BITS'd1524248801, `RNS_PRIME_BITS'd1017883976},
			'{`RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd1036687035, `RNS_PRIME_BITS'd1670803944, `RNS_PRIME_BITS'd700651305, `RNS_PRIME_BITS'd26918801, `RNS_PRIME_BITS'd586065680, `RNS_PRIME_BITS'd1087089814, `RNS_PRIME_BITS'd925328492, `RNS_PRIME_BITS'd754764174, `RNS_PRIME_BITS'd1681243620, `RNS_PRIME_BITS'd207195504},
			'{`RNS_PRIME_BITS'd151, `RNS_PRIME_BITS'd1832917086, `RNS_PRIME_BITS'd797484415, `RNS_PRIME_BITS'd1460028445, `RNS_PRIME_BITS'd215163515, `RNS_PRIME_BITS'd1893508332, `RNS_PRIME_BITS'd826169757, `RNS_PRIME_BITS'd916623069, `RNS_PRIME_BITS'd1118874874, `RNS_PRIME_BITS'd184028124, `RNS_PRIME_BITS'd537079614},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd2078851518, `RNS_PRIME_BITS'd1917046205, `RNS_PRIME_BITS'd1648335652, `RNS_PRIME_BITS'd802596532, `RNS_PRIME_BITS'd1430603199, `RNS_PRIME_BITS'd825058651, `RNS_PRIME_BITS'd1092947588, `RNS_PRIME_BITS'd1162372683, `RNS_PRIME_BITS'd1618224857, `RNS_PRIME_BITS'd505226246},
			'{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd924570036, `RNS_PRIME_BITS'd2120295725, `RNS_PRIME_BITS'd1717858675, `RNS_PRIME_BITS'd1541315518, `RNS_PRIME_BITS'd1383324291, `RNS_PRIME_BITS'd1671357596, `RNS_PRIME_BITS'd628415182, `RNS_PRIME_BITS'd1399526344, `RNS_PRIME_BITS'd2111341219, `RNS_PRIME_BITS'd1876039717},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1522605116, `RNS_PRIME_BITS'd1848997174, `RNS_PRIME_BITS'd1951270127, `RNS_PRIME_BITS'd494520681, `RNS_PRIME_BITS'd1087671684, `RNS_PRIME_BITS'd42778303, `RNS_PRIME_BITS'd1764522565, `RNS_PRIME_BITS'd709852686, `RNS_PRIME_BITS'd1646127238, `RNS_PRIME_BITS'd1800470972},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1945512785, `RNS_PRIME_BITS'd2090804285, `RNS_PRIME_BITS'd1359796239, `RNS_PRIME_BITS'd1042527149, `RNS_PRIME_BITS'd1249094217, `RNS_PRIME_BITS'd576547451, `RNS_PRIME_BITS'd1583629807, `RNS_PRIME_BITS'd1759815402, `RNS_PRIME_BITS'd1904289064, `RNS_PRIME_BITS'd1420160441},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd828294124, `RNS_PRIME_BITS'd802650402, `RNS_PRIME_BITS'd1648561603, `RNS_PRIME_BITS'd234166116, `RNS_PRIME_BITS'd197400809, `RNS_PRIME_BITS'd1903120582, `RNS_PRIME_BITS'd642337414, `RNS_PRIME_BITS'd1934884436, `RNS_PRIME_BITS'd345490476, `RNS_PRIME_BITS'd986146703},
			'{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd774033964, `RNS_PRIME_BITS'd1853787389, `RNS_PRIME_BITS'd1034200850, `RNS_PRIME_BITS'd2003965926, `RNS_PRIME_BITS'd70638059, `RNS_PRIME_BITS'd722824034, `RNS_PRIME_BITS'd1095652287, `RNS_PRIME_BITS'd874915222, `RNS_PRIME_BITS'd2116168641, `RNS_PRIME_BITS'd593671560},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1989762631, `RNS_PRIME_BITS'd926777446, `RNS_PRIME_BITS'd924424222, `RNS_PRIME_BITS'd917510226, `RNS_PRIME_BITS'd108938286, `RNS_PRIME_BITS'd68429361, `RNS_PRIME_BITS'd369886156, `RNS_PRIME_BITS'd682522457, `RNS_PRIME_BITS'd576194945, `RNS_PRIME_BITS'd756290639},
			'{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd900058570, `RNS_PRIME_BITS'd2049655831, `RNS_PRIME_BITS'd549533888, `RNS_PRIME_BITS'd1352964446, `RNS_PRIME_BITS'd1660536834, `RNS_PRIME_BITS'd589288740, `RNS_PRIME_BITS'd531939731, `RNS_PRIME_BITS'd97187497, `RNS_PRIME_BITS'd137299689, `RNS_PRIME_BITS'd1460385311},
			'{`RNS_PRIME_BITS'd156, `RNS_PRIME_BITS'd614467045, `RNS_PRIME_BITS'd1467150196, `RNS_PRIME_BITS'd409453136, `RNS_PRIME_BITS'd430991850, `RNS_PRIME_BITS'd1637818519, `RNS_PRIME_BITS'd1578470715, `RNS_PRIME_BITS'd1683527210, `RNS_PRIME_BITS'd2044955390, `RNS_PRIME_BITS'd1991178869, `RNS_PRIME_BITS'd1282166198},
			'{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd1697668479, `RNS_PRIME_BITS'd1838113925, `RNS_PRIME_BITS'd189158759, `RNS_PRIME_BITS'd788672247, `RNS_PRIME_BITS'd1036320379, `RNS_PRIME_BITS'd665417193, `RNS_PRIME_BITS'd2012864420, `RNS_PRIME_BITS'd1336641007, `RNS_PRIME_BITS'd991058596, `RNS_PRIME_BITS'd127674721},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd1408000316, `RNS_PRIME_BITS'd938536028, `RNS_PRIME_BITS'd1885008653, `RNS_PRIME_BITS'd1352424225, `RNS_PRIME_BITS'd1001621347, `RNS_PRIME_BITS'd204991059, `RNS_PRIME_BITS'd2077001472, `RNS_PRIME_BITS'd236586893, `RNS_PRIME_BITS'd33364519, `RNS_PRIME_BITS'd623856161},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd553862152, `RNS_PRIME_BITS'd155655288, `RNS_PRIME_BITS'd436509812, `RNS_PRIME_BITS'd2094287047, `RNS_PRIME_BITS'd37110479, `RNS_PRIME_BITS'd1373801345, `RNS_PRIME_BITS'd1596098214, `RNS_PRIME_BITS'd736478187, `RNS_PRIME_BITS'd1600443514, `RNS_PRIME_BITS'd1328844776},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd1526513425, `RNS_PRIME_BITS'd2107092954, `RNS_PRIME_BITS'd1733932873, `RNS_PRIME_BITS'd894293400, `RNS_PRIME_BITS'd858879269, `RNS_PRIME_BITS'd166422522, `RNS_PRIME_BITS'd1633913716, `RNS_PRIME_BITS'd1564310417, `RNS_PRIME_BITS'd1739949914, `RNS_PRIME_BITS'd1462167084},
			'{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd1937373608, `RNS_PRIME_BITS'd1072497198, `RNS_PRIME_BITS'd780367099, `RNS_PRIME_BITS'd644429847, `RNS_PRIME_BITS'd651284630, `RNS_PRIME_BITS'd2007872484, `RNS_PRIME_BITS'd664828861, `RNS_PRIME_BITS'd1850282023, `RNS_PRIME_BITS'd661692327, `RNS_PRIME_BITS'd269170542},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd1959357099, `RNS_PRIME_BITS'd950283428, `RNS_PRIME_BITS'd809388721, `RNS_PRIME_BITS'd433974139, `RNS_PRIME_BITS'd1522020410, `RNS_PRIME_BITS'd2020713986, `RNS_PRIME_BITS'd280681878, `RNS_PRIME_BITS'd673228011, `RNS_PRIME_BITS'd2136124212, `RNS_PRIME_BITS'd169483342},
			'{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd10065796, `RNS_PRIME_BITS'd1763431582, `RNS_PRIME_BITS'd1501660343, `RNS_PRIME_BITS'd55855173, `RNS_PRIME_BITS'd1682881588, `RNS_PRIME_BITS'd1303734102, `RNS_PRIME_BITS'd309079992, `RNS_PRIME_BITS'd20143732, `RNS_PRIME_BITS'd1024097300, `RNS_PRIME_BITS'd551406687},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd95534702, `RNS_PRIME_BITS'd1123443552, `RNS_PRIME_BITS'd922259314, `RNS_PRIME_BITS'd1300049469, `RNS_PRIME_BITS'd699418356, `RNS_PRIME_BITS'd1408649948, `RNS_PRIME_BITS'd612087915, `RNS_PRIME_BITS'd1568613164, `RNS_PRIME_BITS'd730048134, `RNS_PRIME_BITS'd1070767751},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1767129584, `RNS_PRIME_BITS'd1299222566, `RNS_PRIME_BITS'd924168161, `RNS_PRIME_BITS'd501752132, `RNS_PRIME_BITS'd939209593, `RNS_PRIME_BITS'd448557300, `RNS_PRIME_BITS'd1016780559, `RNS_PRIME_BITS'd1669199544, `RNS_PRIME_BITS'd2020991252, `RNS_PRIME_BITS'd842714821},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd844473131, `RNS_PRIME_BITS'd553337094, `RNS_PRIME_BITS'd529401120, `RNS_PRIME_BITS'd787400088, `RNS_PRIME_BITS'd2098885882, `RNS_PRIME_BITS'd21834480, `RNS_PRIME_BITS'd132933, `RNS_PRIME_BITS'd1986703582, `RNS_PRIME_BITS'd664929311, `RNS_PRIME_BITS'd1706796478},
			'{`RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd1640063271, `RNS_PRIME_BITS'd1860771052, `RNS_PRIME_BITS'd833777990, `RNS_PRIME_BITS'd490152901, `RNS_PRIME_BITS'd1997034852, `RNS_PRIME_BITS'd1805239800, `RNS_PRIME_BITS'd2033332974, `RNS_PRIME_BITS'd1456427129, `RNS_PRIME_BITS'd478701145, `RNS_PRIME_BITS'd801911286},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd1308180011, `RNS_PRIME_BITS'd735084563, `RNS_PRIME_BITS'd1329547201, `RNS_PRIME_BITS'd821721125, `RNS_PRIME_BITS'd138231851, `RNS_PRIME_BITS'd892360492, `RNS_PRIME_BITS'd1484336147, `RNS_PRIME_BITS'd249176400, `RNS_PRIME_BITS'd2074587080, `RNS_PRIME_BITS'd1482841647},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd1497855394, `RNS_PRIME_BITS'd1942273652, `RNS_PRIME_BITS'd724532963, `RNS_PRIME_BITS'd901967230, `RNS_PRIME_BITS'd1392289554, `RNS_PRIME_BITS'd1029947084, `RNS_PRIME_BITS'd1014455886, `RNS_PRIME_BITS'd1505151617, `RNS_PRIME_BITS'd1437173336, `RNS_PRIME_BITS'd280692357},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd416804320, `RNS_PRIME_BITS'd1177683841, `RNS_PRIME_BITS'd742986795, `RNS_PRIME_BITS'd1743136356, `RNS_PRIME_BITS'd1564759358, `RNS_PRIME_BITS'd280471959, `RNS_PRIME_BITS'd1039640051, `RNS_PRIME_BITS'd14550967, `RNS_PRIME_BITS'd576995966, `RNS_PRIME_BITS'd1785629487},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1288144363, `RNS_PRIME_BITS'd1281603594, `RNS_PRIME_BITS'd2071198473, `RNS_PRIME_BITS'd1908089657, `RNS_PRIME_BITS'd302611111, `RNS_PRIME_BITS'd924399381, `RNS_PRIME_BITS'd724804413, `RNS_PRIME_BITS'd1953358574, `RNS_PRIME_BITS'd690463787, `RNS_PRIME_BITS'd1464689878},
			'{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd956116996, `RNS_PRIME_BITS'd684747443, `RNS_PRIME_BITS'd1412426776, `RNS_PRIME_BITS'd8357172, `RNS_PRIME_BITS'd618260026, `RNS_PRIME_BITS'd142597389, `RNS_PRIME_BITS'd895167180, `RNS_PRIME_BITS'd1443130654, `RNS_PRIME_BITS'd66475800, `RNS_PRIME_BITS'd1711047663},
			'{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd1649696949, `RNS_PRIME_BITS'd1464510865, `RNS_PRIME_BITS'd1206309906, `RNS_PRIME_BITS'd1746424778, `RNS_PRIME_BITS'd1994753370, `RNS_PRIME_BITS'd59942719, `RNS_PRIME_BITS'd558509959, `RNS_PRIME_BITS'd1565938580, `RNS_PRIME_BITS'd330950088, `RNS_PRIME_BITS'd1336355439},
			'{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd1820359959, `RNS_PRIME_BITS'd1180814713, `RNS_PRIME_BITS'd1743628342, `RNS_PRIME_BITS'd421534736, `RNS_PRIME_BITS'd1150168763, `RNS_PRIME_BITS'd1266369661, `RNS_PRIME_BITS'd2076760559, `RNS_PRIME_BITS'd1000841432, `RNS_PRIME_BITS'd335583260, `RNS_PRIME_BITS'd929426088},
			'{`RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd758900630, `RNS_PRIME_BITS'd673236382, `RNS_PRIME_BITS'd346682446, `RNS_PRIME_BITS'd696468798, `RNS_PRIME_BITS'd294060537, `RNS_PRIME_BITS'd1458044052, `RNS_PRIME_BITS'd1372476949, `RNS_PRIME_BITS'd1249841786, `RNS_PRIME_BITS'd443380456, `RNS_PRIME_BITS'd98314169},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1287307662, `RNS_PRIME_BITS'd1973595280, `RNS_PRIME_BITS'd175265562, `RNS_PRIME_BITS'd2067234556, `RNS_PRIME_BITS'd1234926776, `RNS_PRIME_BITS'd283840506, `RNS_PRIME_BITS'd882254174, `RNS_PRIME_BITS'd1859536826, `RNS_PRIME_BITS'd695995556, `RNS_PRIME_BITS'd1679292023},
			'{`RNS_PRIME_BITS'd169, `RNS_PRIME_BITS'd429039396, `RNS_PRIME_BITS'd818944881, `RNS_PRIME_BITS'd868918149, `RNS_PRIME_BITS'd1505651808, `RNS_PRIME_BITS'd2137491613, `RNS_PRIME_BITS'd185431750, `RNS_PRIME_BITS'd985768460, `RNS_PRIME_BITS'd326774881, `RNS_PRIME_BITS'd1937138814, `RNS_PRIME_BITS'd48653958},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd999033149, `RNS_PRIME_BITS'd1891695094, `RNS_PRIME_BITS'd1370889966, `RNS_PRIME_BITS'd592767796, `RNS_PRIME_BITS'd1993577447, `RNS_PRIME_BITS'd1430559940, `RNS_PRIME_BITS'd2081084747, `RNS_PRIME_BITS'd490567660, `RNS_PRIME_BITS'd1090546565, `RNS_PRIME_BITS'd858163832},
			'{`RNS_PRIME_BITS'd196, `RNS_PRIME_BITS'd1386979332, `RNS_PRIME_BITS'd1121970187, `RNS_PRIME_BITS'd232318749, `RNS_PRIME_BITS'd672623745, `RNS_PRIME_BITS'd1733057332, `RNS_PRIME_BITS'd1373999916, `RNS_PRIME_BITS'd1437233917, `RNS_PRIME_BITS'd574670363, `RNS_PRIME_BITS'd680467917, `RNS_PRIME_BITS'd1944373885},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd1779724213, `RNS_PRIME_BITS'd2101086503, `RNS_PRIME_BITS'd379592967, `RNS_PRIME_BITS'd2089704760, `RNS_PRIME_BITS'd2032096005, `RNS_PRIME_BITS'd1166156876, `RNS_PRIME_BITS'd2098766330, `RNS_PRIME_BITS'd1957490628, `RNS_PRIME_BITS'd1437896994, `RNS_PRIME_BITS'd1195203553},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd1307574237, `RNS_PRIME_BITS'd634066391, `RNS_PRIME_BITS'd765851082, `RNS_PRIME_BITS'd1790367302, `RNS_PRIME_BITS'd1630996790, `RNS_PRIME_BITS'd290130221, `RNS_PRIME_BITS'd15991371, `RNS_PRIME_BITS'd1166213289, `RNS_PRIME_BITS'd1460870024, `RNS_PRIME_BITS'd1092038724}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd1460001394, `RNS_PRIME_BITS'd315111235, `RNS_PRIME_BITS'd1770527196, `RNS_PRIME_BITS'd1654653288, `RNS_PRIME_BITS'd1964852308, `RNS_PRIME_BITS'd1658430858, `RNS_PRIME_BITS'd131163702, `RNS_PRIME_BITS'd287182049, `RNS_PRIME_BITS'd1930009758, `RNS_PRIME_BITS'd743552137},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1316075784, `RNS_PRIME_BITS'd657559923, `RNS_PRIME_BITS'd2139882512, `RNS_PRIME_BITS'd700195685, `RNS_PRIME_BITS'd874424013, `RNS_PRIME_BITS'd701669091, `RNS_PRIME_BITS'd1479657245, `RNS_PRIME_BITS'd470523888, `RNS_PRIME_BITS'd920635718, `RNS_PRIME_BITS'd785438018},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd525546596, `RNS_PRIME_BITS'd268111859, `RNS_PRIME_BITS'd1570610927, `RNS_PRIME_BITS'd472257421, `RNS_PRIME_BITS'd1350708573, `RNS_PRIME_BITS'd1685219791, `RNS_PRIME_BITS'd1813662886, `RNS_PRIME_BITS'd273109519, `RNS_PRIME_BITS'd1217984333, `RNS_PRIME_BITS'd1745945767},
			'{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd491708291, `RNS_PRIME_BITS'd1224216088, `RNS_PRIME_BITS'd800568893, `RNS_PRIME_BITS'd1287059478, `RNS_PRIME_BITS'd1530154018, `RNS_PRIME_BITS'd519356292, `RNS_PRIME_BITS'd923491777, `RNS_PRIME_BITS'd1722839936, `RNS_PRIME_BITS'd1691135635, `RNS_PRIME_BITS'd593404540},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1231033388, `RNS_PRIME_BITS'd1767872324, `RNS_PRIME_BITS'd1493140125, `RNS_PRIME_BITS'd1846978952, `RNS_PRIME_BITS'd718482450, `RNS_PRIME_BITS'd548467401, `RNS_PRIME_BITS'd2028897087, `RNS_PRIME_BITS'd1628791628, `RNS_PRIME_BITS'd1855185269, `RNS_PRIME_BITS'd15225243},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1439054782, `RNS_PRIME_BITS'd766360626, `RNS_PRIME_BITS'd1968342993, `RNS_PRIME_BITS'd2043489572, `RNS_PRIME_BITS'd412325835, `RNS_PRIME_BITS'd171387828, `RNS_PRIME_BITS'd1817062841, `RNS_PRIME_BITS'd197715351, `RNS_PRIME_BITS'd1696069699, `RNS_PRIME_BITS'd1057709687},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd422060688, `RNS_PRIME_BITS'd1316645531, `RNS_PRIME_BITS'd578543145, `RNS_PRIME_BITS'd813164106, `RNS_PRIME_BITS'd1506514821, `RNS_PRIME_BITS'd786602513, `RNS_PRIME_BITS'd19007350, `RNS_PRIME_BITS'd1328635300, `RNS_PRIME_BITS'd1349511362, `RNS_PRIME_BITS'd458324330},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd1461014953, `RNS_PRIME_BITS'd2057415366, `RNS_PRIME_BITS'd1656034993, `RNS_PRIME_BITS'd919707778, `RNS_PRIME_BITS'd822591332, `RNS_PRIME_BITS'd1359550384, `RNS_PRIME_BITS'd877125005, `RNS_PRIME_BITS'd957296449, `RNS_PRIME_BITS'd658704943, `RNS_PRIME_BITS'd766136866},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1993180374, `RNS_PRIME_BITS'd1175841003, `RNS_PRIME_BITS'd662999838, `RNS_PRIME_BITS'd595382293, `RNS_PRIME_BITS'd1766082488, `RNS_PRIME_BITS'd863807213, `RNS_PRIME_BITS'd1244961774, `RNS_PRIME_BITS'd1325264013, `RNS_PRIME_BITS'd1832509498, `RNS_PRIME_BITS'd122188539},
			'{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd1795197597, `RNS_PRIME_BITS'd1541428075, `RNS_PRIME_BITS'd825392396, `RNS_PRIME_BITS'd1945101182, `RNS_PRIME_BITS'd2098661277, `RNS_PRIME_BITS'd307290991, `RNS_PRIME_BITS'd204538861, `RNS_PRIME_BITS'd1552032846, `RNS_PRIME_BITS'd1658765590, `RNS_PRIME_BITS'd777961599},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1920080172, `RNS_PRIME_BITS'd2023028706, `RNS_PRIME_BITS'd537323821, `RNS_PRIME_BITS'd929501402, `RNS_PRIME_BITS'd1400135286, `RNS_PRIME_BITS'd197670302, `RNS_PRIME_BITS'd1486503342, `RNS_PRIME_BITS'd2073170930, `RNS_PRIME_BITS'd1781620271, `RNS_PRIME_BITS'd603845659},
			'{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd92798718, `RNS_PRIME_BITS'd353896536, `RNS_PRIME_BITS'd653077770, `RNS_PRIME_BITS'd1219656882, `RNS_PRIME_BITS'd82294942, `RNS_PRIME_BITS'd499521962, `RNS_PRIME_BITS'd1370038664, `RNS_PRIME_BITS'd1648205026, `RNS_PRIME_BITS'd1492362339, `RNS_PRIME_BITS'd294308935},
			'{`RNS_PRIME_BITS'd127, `RNS_PRIME_BITS'd55826711, `RNS_PRIME_BITS'd863035292, `RNS_PRIME_BITS'd355436969, `RNS_PRIME_BITS'd1712110623, `RNS_PRIME_BITS'd1182417624, `RNS_PRIME_BITS'd930811885, `RNS_PRIME_BITS'd767935667, `RNS_PRIME_BITS'd1265121556, `RNS_PRIME_BITS'd770081760, `RNS_PRIME_BITS'd1644159064},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd531783944, `RNS_PRIME_BITS'd1395008889, `RNS_PRIME_BITS'd1921838443, `RNS_PRIME_BITS'd450742121, `RNS_PRIME_BITS'd1624054564, `RNS_PRIME_BITS'd124231665, `RNS_PRIME_BITS'd1491338779, `RNS_PRIME_BITS'd1087003959, `RNS_PRIME_BITS'd394712780, `RNS_PRIME_BITS'd1818106137},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd1115029187, `RNS_PRIME_BITS'd1865758534, `RNS_PRIME_BITS'd1040290429, `RNS_PRIME_BITS'd440868770, `RNS_PRIME_BITS'd1754116729, `RNS_PRIME_BITS'd16426510, `RNS_PRIME_BITS'd45208685, `RNS_PRIME_BITS'd1809260565, `RNS_PRIME_BITS'd573136611, `RNS_PRIME_BITS'd1930048231},
			'{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd30484207, `RNS_PRIME_BITS'd544136084, `RNS_PRIME_BITS'd1249838004, `RNS_PRIME_BITS'd2051416705, `RNS_PRIME_BITS'd1286129451, `RNS_PRIME_BITS'd200693587, `RNS_PRIME_BITS'd1261695839, `RNS_PRIME_BITS'd1906500233, `RNS_PRIME_BITS'd1309945706, `RNS_PRIME_BITS'd1158926112},
			'{`RNS_PRIME_BITS'd63, `RNS_PRIME_BITS'd862269045, `RNS_PRIME_BITS'd441535876, `RNS_PRIME_BITS'd890269683, `RNS_PRIME_BITS'd637194158, `RNS_PRIME_BITS'd361856850, `RNS_PRIME_BITS'd2073245316, `RNS_PRIME_BITS'd2056622534, `RNS_PRIME_BITS'd1188063834, `RNS_PRIME_BITS'd90943457, `RNS_PRIME_BITS'd109452174},
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd1936406680, `RNS_PRIME_BITS'd685813054, `RNS_PRIME_BITS'd1435309695, `RNS_PRIME_BITS'd1597636721, `RNS_PRIME_BITS'd581199048, `RNS_PRIME_BITS'd189982621, `RNS_PRIME_BITS'd1206186630, `RNS_PRIME_BITS'd1855175424, `RNS_PRIME_BITS'd1066328376, `RNS_PRIME_BITS'd1644323983},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd416422674, `RNS_PRIME_BITS'd40079743, `RNS_PRIME_BITS'd1424231425, `RNS_PRIME_BITS'd95461318, `RNS_PRIME_BITS'd1383660014, `RNS_PRIME_BITS'd1499895471, `RNS_PRIME_BITS'd82454295, `RNS_PRIME_BITS'd153531259, `RNS_PRIME_BITS'd217942645, `RNS_PRIME_BITS'd216764268},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1403220007, `RNS_PRIME_BITS'd1312232701, `RNS_PRIME_BITS'd214280685, `RNS_PRIME_BITS'd218300651, `RNS_PRIME_BITS'd801795142, `RNS_PRIME_BITS'd1921378331, `RNS_PRIME_BITS'd898429609, `RNS_PRIME_BITS'd652911729, `RNS_PRIME_BITS'd1562248329, `RNS_PRIME_BITS'd1514470789},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd1653228724, `RNS_PRIME_BITS'd680518544, `RNS_PRIME_BITS'd1555908402, `RNS_PRIME_BITS'd1730867477, `RNS_PRIME_BITS'd125396276, `RNS_PRIME_BITS'd626235030, `RNS_PRIME_BITS'd1559305718, `RNS_PRIME_BITS'd65267805, `RNS_PRIME_BITS'd713509644, `RNS_PRIME_BITS'd749666972},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1904819856, `RNS_PRIME_BITS'd1598097705, `RNS_PRIME_BITS'd849568577, `RNS_PRIME_BITS'd1623731489, `RNS_PRIME_BITS'd1092573723, `RNS_PRIME_BITS'd1183341120, `RNS_PRIME_BITS'd517243304, `RNS_PRIME_BITS'd833203219, `RNS_PRIME_BITS'd403924833, `RNS_PRIME_BITS'd601872792},
			'{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd776592907, `RNS_PRIME_BITS'd1299747487, `RNS_PRIME_BITS'd1489051909, `RNS_PRIME_BITS'd488915692, `RNS_PRIME_BITS'd943191861, `RNS_PRIME_BITS'd1663719710, `RNS_PRIME_BITS'd651093936, `RNS_PRIME_BITS'd624817483, `RNS_PRIME_BITS'd1198814570, `RNS_PRIME_BITS'd1573982316},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1244631163, `RNS_PRIME_BITS'd507386565, `RNS_PRIME_BITS'd1324826333, `RNS_PRIME_BITS'd1041463192, `RNS_PRIME_BITS'd1351766057, `RNS_PRIME_BITS'd1930784064, `RNS_PRIME_BITS'd2014156290, `RNS_PRIME_BITS'd296937981, `RNS_PRIME_BITS'd768847601, `RNS_PRIME_BITS'd88691188},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd1593249079, `RNS_PRIME_BITS'd460997180, `RNS_PRIME_BITS'd1286763700, `RNS_PRIME_BITS'd878571718, `RNS_PRIME_BITS'd1456909119, `RNS_PRIME_BITS'd801219748, `RNS_PRIME_BITS'd1574359378, `RNS_PRIME_BITS'd1112391338, `RNS_PRIME_BITS'd979008445, `RNS_PRIME_BITS'd1516251896},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd1417015336, `RNS_PRIME_BITS'd1631485882, `RNS_PRIME_BITS'd1537188679, `RNS_PRIME_BITS'd32701206, `RNS_PRIME_BITS'd941769400, `RNS_PRIME_BITS'd1979318650, `RNS_PRIME_BITS'd213563633, `RNS_PRIME_BITS'd721109361, `RNS_PRIME_BITS'd1482829175, `RNS_PRIME_BITS'd898927783},
			'{`RNS_PRIME_BITS'd109, `RNS_PRIME_BITS'd338277351, `RNS_PRIME_BITS'd253122682, `RNS_PRIME_BITS'd1959677985, `RNS_PRIME_BITS'd580264481, `RNS_PRIME_BITS'd785440066, `RNS_PRIME_BITS'd1444412439, `RNS_PRIME_BITS'd1123039323, `RNS_PRIME_BITS'd1297770788, `RNS_PRIME_BITS'd1488886017, `RNS_PRIME_BITS'd1101002870},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1471591937, `RNS_PRIME_BITS'd358551347, `RNS_PRIME_BITS'd490798113, `RNS_PRIME_BITS'd1362350796, `RNS_PRIME_BITS'd1275231291, `RNS_PRIME_BITS'd1428111266, `RNS_PRIME_BITS'd745825073, `RNS_PRIME_BITS'd391664885, `RNS_PRIME_BITS'd2019200783, `RNS_PRIME_BITS'd485741706},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd663743728, `RNS_PRIME_BITS'd108360531, `RNS_PRIME_BITS'd1184127399, `RNS_PRIME_BITS'd2124915455, `RNS_PRIME_BITS'd2034502074, `RNS_PRIME_BITS'd802773450, `RNS_PRIME_BITS'd1339693456, `RNS_PRIME_BITS'd1865394147, `RNS_PRIME_BITS'd649167475, `RNS_PRIME_BITS'd1612701620},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd2053407303, `RNS_PRIME_BITS'd1443733517, `RNS_PRIME_BITS'd1860911715, `RNS_PRIME_BITS'd2055727854, `RNS_PRIME_BITS'd477942089, `RNS_PRIME_BITS'd1447822413, `RNS_PRIME_BITS'd1725228064, `RNS_PRIME_BITS'd117282573, `RNS_PRIME_BITS'd1444186545, `RNS_PRIME_BITS'd584869042},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd1625198248, `RNS_PRIME_BITS'd1049015575, `RNS_PRIME_BITS'd680830404, `RNS_PRIME_BITS'd1955717997, `RNS_PRIME_BITS'd259494093, `RNS_PRIME_BITS'd1325306881, `RNS_PRIME_BITS'd1040401027, `RNS_PRIME_BITS'd2102621093, `RNS_PRIME_BITS'd2051355854, `RNS_PRIME_BITS'd1600102097},
			'{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd789713422, `RNS_PRIME_BITS'd122271488, `RNS_PRIME_BITS'd1894633858, `RNS_PRIME_BITS'd2140517067, `RNS_PRIME_BITS'd144235241, `RNS_PRIME_BITS'd1159473000, `RNS_PRIME_BITS'd1348625768, `RNS_PRIME_BITS'd1372950652, `RNS_PRIME_BITS'd13626774, `RNS_PRIME_BITS'd696775752},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd313730943, `RNS_PRIME_BITS'd1159891251, `RNS_PRIME_BITS'd906840473, `RNS_PRIME_BITS'd195401283, `RNS_PRIME_BITS'd265515258, `RNS_PRIME_BITS'd1390128889, `RNS_PRIME_BITS'd693858566, `RNS_PRIME_BITS'd1266861147, `RNS_PRIME_BITS'd1774732263, `RNS_PRIME_BITS'd1668560711},
			'{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd833223617, `RNS_PRIME_BITS'd1355973413, `RNS_PRIME_BITS'd1105174380, `RNS_PRIME_BITS'd1143759897, `RNS_PRIME_BITS'd1631841256, `RNS_PRIME_BITS'd2109298418, `RNS_PRIME_BITS'd672141786, `RNS_PRIME_BITS'd918930569, `RNS_PRIME_BITS'd759837144, `RNS_PRIME_BITS'd796872113},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd771783873, `RNS_PRIME_BITS'd1654959120, `RNS_PRIME_BITS'd1631857160, `RNS_PRIME_BITS'd865139934, `RNS_PRIME_BITS'd549737007, `RNS_PRIME_BITS'd1924077826, `RNS_PRIME_BITS'd693065353, `RNS_PRIME_BITS'd110684187, `RNS_PRIME_BITS'd1679802001, `RNS_PRIME_BITS'd698125501},
			'{`RNS_PRIME_BITS'd98, `RNS_PRIME_BITS'd1319572831, `RNS_PRIME_BITS'd330285973, `RNS_PRIME_BITS'd1979898810, `RNS_PRIME_BITS'd715202002, `RNS_PRIME_BITS'd1211264719, `RNS_PRIME_BITS'd328815584, `RNS_PRIME_BITS'd2132787869, `RNS_PRIME_BITS'd2136645431, `RNS_PRIME_BITS'd213269982, `RNS_PRIME_BITS'd691187451},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd2074017676, `RNS_PRIME_BITS'd780155636, `RNS_PRIME_BITS'd992274248, `RNS_PRIME_BITS'd1114943335, `RNS_PRIME_BITS'd1730678341, `RNS_PRIME_BITS'd1928872426, `RNS_PRIME_BITS'd2104726958, `RNS_PRIME_BITS'd1931579267, `RNS_PRIME_BITS'd1317796865, `RNS_PRIME_BITS'd547015746},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd214683641, `RNS_PRIME_BITS'd2038882056, `RNS_PRIME_BITS'd360235563, `RNS_PRIME_BITS'd378231538, `RNS_PRIME_BITS'd1758307065, `RNS_PRIME_BITS'd2145229888, `RNS_PRIME_BITS'd1149108141, `RNS_PRIME_BITS'd1572023709, `RNS_PRIME_BITS'd1641064693, `RNS_PRIME_BITS'd296200014},
			'{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd1592652879, `RNS_PRIME_BITS'd1487707660, `RNS_PRIME_BITS'd1398370530, `RNS_PRIME_BITS'd1970352333, `RNS_PRIME_BITS'd1374971744, `RNS_PRIME_BITS'd245490169, `RNS_PRIME_BITS'd1330256041, `RNS_PRIME_BITS'd436619231, `RNS_PRIME_BITS'd802469311, `RNS_PRIME_BITS'd1272768159},
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd1143578163, `RNS_PRIME_BITS'd1833212924, `RNS_PRIME_BITS'd1291685599, `RNS_PRIME_BITS'd1868008168, `RNS_PRIME_BITS'd1622837818, `RNS_PRIME_BITS'd1956160541, `RNS_PRIME_BITS'd891379127, `RNS_PRIME_BITS'd1725807806, `RNS_PRIME_BITS'd1420238, `RNS_PRIME_BITS'd881911573},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd402943221, `RNS_PRIME_BITS'd1630908627, `RNS_PRIME_BITS'd2002846945, `RNS_PRIME_BITS'd737032397, `RNS_PRIME_BITS'd1233887882, `RNS_PRIME_BITS'd1888970782, `RNS_PRIME_BITS'd1797017821, `RNS_PRIME_BITS'd1555418875, `RNS_PRIME_BITS'd2091741324, `RNS_PRIME_BITS'd480373675},
			'{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd1553191577, `RNS_PRIME_BITS'd870296125, `RNS_PRIME_BITS'd957249438, `RNS_PRIME_BITS'd660190781, `RNS_PRIME_BITS'd1079677161, `RNS_PRIME_BITS'd1680792516, `RNS_PRIME_BITS'd1585346916, `RNS_PRIME_BITS'd1414742800, `RNS_PRIME_BITS'd1516430248, `RNS_PRIME_BITS'd888004993},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd499437665, `RNS_PRIME_BITS'd458956142, `RNS_PRIME_BITS'd272977150, `RNS_PRIME_BITS'd974373343, `RNS_PRIME_BITS'd81013831, `RNS_PRIME_BITS'd1887419821, `RNS_PRIME_BITS'd18205249, `RNS_PRIME_BITS'd224211959, `RNS_PRIME_BITS'd1872659191, `RNS_PRIME_BITS'd1750097568},
			'{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd1666667315, `RNS_PRIME_BITS'd2036691988, `RNS_PRIME_BITS'd597291115, `RNS_PRIME_BITS'd507177022, `RNS_PRIME_BITS'd213424747, `RNS_PRIME_BITS'd140559356, `RNS_PRIME_BITS'd1952513516, `RNS_PRIME_BITS'd1403398798, `RNS_PRIME_BITS'd228664362, `RNS_PRIME_BITS'd1537596429},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd170935425, `RNS_PRIME_BITS'd1412248367, `RNS_PRIME_BITS'd972201676, `RNS_PRIME_BITS'd307697355, `RNS_PRIME_BITS'd651468218, `RNS_PRIME_BITS'd1466547929, `RNS_PRIME_BITS'd244363024, `RNS_PRIME_BITS'd1903510152, `RNS_PRIME_BITS'd102805179, `RNS_PRIME_BITS'd1071560693},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd681202570, `RNS_PRIME_BITS'd77125639, `RNS_PRIME_BITS'd1381754470, `RNS_PRIME_BITS'd418876234, `RNS_PRIME_BITS'd1466338187, `RNS_PRIME_BITS'd955703003, `RNS_PRIME_BITS'd22929632, `RNS_PRIME_BITS'd1871795658, `RNS_PRIME_BITS'd435882375, `RNS_PRIME_BITS'd848205153},
			'{`RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd371348061, `RNS_PRIME_BITS'd295472678, `RNS_PRIME_BITS'd1726142647, `RNS_PRIME_BITS'd1023242696, `RNS_PRIME_BITS'd94368525, `RNS_PRIME_BITS'd2035670113, `RNS_PRIME_BITS'd30194085, `RNS_PRIME_BITS'd1880469106, `RNS_PRIME_BITS'd718575038, `RNS_PRIME_BITS'd1802660768},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd543939467, `RNS_PRIME_BITS'd1323866406, `RNS_PRIME_BITS'd1043422204, `RNS_PRIME_BITS'd133101628, `RNS_PRIME_BITS'd1416487554, `RNS_PRIME_BITS'd424287337, `RNS_PRIME_BITS'd1279431832, `RNS_PRIME_BITS'd1285327152, `RNS_PRIME_BITS'd2013342430, `RNS_PRIME_BITS'd874913289},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1326983414, `RNS_PRIME_BITS'd1064013187, `RNS_PRIME_BITS'd1572843779, `RNS_PRIME_BITS'd1677562397, `RNS_PRIME_BITS'd675940510, `RNS_PRIME_BITS'd290614321, `RNS_PRIME_BITS'd1520932301, `RNS_PRIME_BITS'd391136134, `RNS_PRIME_BITS'd2049041629, `RNS_PRIME_BITS'd1763270999},
			'{`RNS_PRIME_BITS'd54, `RNS_PRIME_BITS'd236684090, `RNS_PRIME_BITS'd834794840, `RNS_PRIME_BITS'd842239864, `RNS_PRIME_BITS'd819244379, `RNS_PRIME_BITS'd1702616229, `RNS_PRIME_BITS'd271702650, `RNS_PRIME_BITS'd1036554475, `RNS_PRIME_BITS'd445722873, `RNS_PRIME_BITS'd1921855870, `RNS_PRIME_BITS'd1877204802},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd874930695, `RNS_PRIME_BITS'd905507326, `RNS_PRIME_BITS'd145039391, `RNS_PRIME_BITS'd1386090509, `RNS_PRIME_BITS'd2121510301, `RNS_PRIME_BITS'd109085205, `RNS_PRIME_BITS'd710521979, `RNS_PRIME_BITS'd4702437, `RNS_PRIME_BITS'd760442202, `RNS_PRIME_BITS'd241809229},
			'{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd1956922989, `RNS_PRIME_BITS'd885086663, `RNS_PRIME_BITS'd1496010882, `RNS_PRIME_BITS'd870280648, `RNS_PRIME_BITS'd1446654199, `RNS_PRIME_BITS'd1872883954, `RNS_PRIME_BITS'd1519143761, `RNS_PRIME_BITS'd961624685, `RNS_PRIME_BITS'd1967959676, `RNS_PRIME_BITS'd1373556750},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1338232044, `RNS_PRIME_BITS'd1322475571, `RNS_PRIME_BITS'd2059570337, `RNS_PRIME_BITS'd1943495341, `RNS_PRIME_BITS'd822335282, `RNS_PRIME_BITS'd1628701385, `RNS_PRIME_BITS'd807026028, `RNS_PRIME_BITS'd1259810574, `RNS_PRIME_BITS'd1961811113, `RNS_PRIME_BITS'd783603009},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd991602813, `RNS_PRIME_BITS'd353965818, `RNS_PRIME_BITS'd1574054566, `RNS_PRIME_BITS'd812830933, `RNS_PRIME_BITS'd1477655043, `RNS_PRIME_BITS'd472001571, `RNS_PRIME_BITS'd1423892519, `RNS_PRIME_BITS'd1351484672, `RNS_PRIME_BITS'd762931885, `RNS_PRIME_BITS'd1299470103},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1266272703, `RNS_PRIME_BITS'd1696724783, `RNS_PRIME_BITS'd1487824757, `RNS_PRIME_BITS'd168853514, `RNS_PRIME_BITS'd961831592, `RNS_PRIME_BITS'd1993028677, `RNS_PRIME_BITS'd841002035, `RNS_PRIME_BITS'd529696984, `RNS_PRIME_BITS'd1601873186, `RNS_PRIME_BITS'd1428705065},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd351347113, `RNS_PRIME_BITS'd1264814131, `RNS_PRIME_BITS'd1471686775, `RNS_PRIME_BITS'd883051146, `RNS_PRIME_BITS'd1454770106, `RNS_PRIME_BITS'd1283105884, `RNS_PRIME_BITS'd610071169, `RNS_PRIME_BITS'd1190020558, `RNS_PRIME_BITS'd434803654, `RNS_PRIME_BITS'd894158025},
			'{`RNS_PRIME_BITS'd188, `RNS_PRIME_BITS'd86779768, `RNS_PRIME_BITS'd1784517486, `RNS_PRIME_BITS'd749053403, `RNS_PRIME_BITS'd1197602312, `RNS_PRIME_BITS'd2009025797, `RNS_PRIME_BITS'd463942571, `RNS_PRIME_BITS'd726577738, `RNS_PRIME_BITS'd1264842667, `RNS_PRIME_BITS'd2118849645, `RNS_PRIME_BITS'd1827858703},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd391227431, `RNS_PRIME_BITS'd1320653066, `RNS_PRIME_BITS'd1849215226, `RNS_PRIME_BITS'd2056850828, `RNS_PRIME_BITS'd270145631, `RNS_PRIME_BITS'd1864427790, `RNS_PRIME_BITS'd1812550297, `RNS_PRIME_BITS'd716012975, `RNS_PRIME_BITS'd1459041617, `RNS_PRIME_BITS'd1574398017},
			'{`RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd1084275408, `RNS_PRIME_BITS'd945147262, `RNS_PRIME_BITS'd1318723069, `RNS_PRIME_BITS'd1332950614, `RNS_PRIME_BITS'd571752776, `RNS_PRIME_BITS'd464857870, `RNS_PRIME_BITS'd1390491869, `RNS_PRIME_BITS'd47344842, `RNS_PRIME_BITS'd1774765877, `RNS_PRIME_BITS'd1621348317},
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd100964001, `RNS_PRIME_BITS'd1107400438, `RNS_PRIME_BITS'd460062096, `RNS_PRIME_BITS'd1308244894, `RNS_PRIME_BITS'd43428190, `RNS_PRIME_BITS'd1145635307, `RNS_PRIME_BITS'd457134637, `RNS_PRIME_BITS'd513494111, `RNS_PRIME_BITS'd264661579, `RNS_PRIME_BITS'd1543430323},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd154494120, `RNS_PRIME_BITS'd1830149911, `RNS_PRIME_BITS'd515188530, `RNS_PRIME_BITS'd1982201173, `RNS_PRIME_BITS'd2050018196, `RNS_PRIME_BITS'd705081211, `RNS_PRIME_BITS'd1981292228, `RNS_PRIME_BITS'd1850370797, `RNS_PRIME_BITS'd228050518, `RNS_PRIME_BITS'd751135560},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd1053371529, `RNS_PRIME_BITS'd543225476, `RNS_PRIME_BITS'd1522036019, `RNS_PRIME_BITS'd1148835249, `RNS_PRIME_BITS'd459147536, `RNS_PRIME_BITS'd585952887, `RNS_PRIME_BITS'd481728279, `RNS_PRIME_BITS'd2059785118, `RNS_PRIME_BITS'd1707530308, `RNS_PRIME_BITS'd665982803},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd1851578048, `RNS_PRIME_BITS'd702920578, `RNS_PRIME_BITS'd1228038389, `RNS_PRIME_BITS'd649971267, `RNS_PRIME_BITS'd322058983, `RNS_PRIME_BITS'd1040280786, `RNS_PRIME_BITS'd171551625, `RNS_PRIME_BITS'd1648588339, `RNS_PRIME_BITS'd1366766655, `RNS_PRIME_BITS'd414382466},
			'{`RNS_PRIME_BITS'd76, `RNS_PRIME_BITS'd577006648, `RNS_PRIME_BITS'd148990400, `RNS_PRIME_BITS'd211641671, `RNS_PRIME_BITS'd959706336, `RNS_PRIME_BITS'd1005740920, `RNS_PRIME_BITS'd271361394, `RNS_PRIME_BITS'd1641194420, `RNS_PRIME_BITS'd1023988028, `RNS_PRIME_BITS'd1132471233, `RNS_PRIME_BITS'd274053565}
		},
		'{
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd1582959541, `RNS_PRIME_BITS'd611154289, `RNS_PRIME_BITS'd895086121, `RNS_PRIME_BITS'd1165253425, `RNS_PRIME_BITS'd1839947582, `RNS_PRIME_BITS'd1004427184, `RNS_PRIME_BITS'd574266707, `RNS_PRIME_BITS'd1852128302, `RNS_PRIME_BITS'd491393687, `RNS_PRIME_BITS'd50960693},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd260740311, `RNS_PRIME_BITS'd79875103, `RNS_PRIME_BITS'd141374794, `RNS_PRIME_BITS'd224085048, `RNS_PRIME_BITS'd1829974560, `RNS_PRIME_BITS'd781744180, `RNS_PRIME_BITS'd1323329435, `RNS_PRIME_BITS'd628886928, `RNS_PRIME_BITS'd1431510646, `RNS_PRIME_BITS'd1250808217},
			'{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd1562013821, `RNS_PRIME_BITS'd761437878, `RNS_PRIME_BITS'd1819814443, `RNS_PRIME_BITS'd1620007936, `RNS_PRIME_BITS'd1169851131, `RNS_PRIME_BITS'd207230025, `RNS_PRIME_BITS'd1170592130, `RNS_PRIME_BITS'd311629980, `RNS_PRIME_BITS'd1034119553, `RNS_PRIME_BITS'd1706224830},
			'{`RNS_PRIME_BITS'd188, `RNS_PRIME_BITS'd1014828462, `RNS_PRIME_BITS'd1814563623, `RNS_PRIME_BITS'd1759580452, `RNS_PRIME_BITS'd1477649288, `RNS_PRIME_BITS'd971991568, `RNS_PRIME_BITS'd2040138734, `RNS_PRIME_BITS'd550407712, `RNS_PRIME_BITS'd1502941429, `RNS_PRIME_BITS'd2003261959, `RNS_PRIME_BITS'd1992814006},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd92950919, `RNS_PRIME_BITS'd1977070716, `RNS_PRIME_BITS'd676964094, `RNS_PRIME_BITS'd521884396, `RNS_PRIME_BITS'd1401714691, `RNS_PRIME_BITS'd974197549, `RNS_PRIME_BITS'd906143825, `RNS_PRIME_BITS'd1757743207, `RNS_PRIME_BITS'd898892247, `RNS_PRIME_BITS'd198127091},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd2070008811, `RNS_PRIME_BITS'd8161822, `RNS_PRIME_BITS'd605698489, `RNS_PRIME_BITS'd566743395, `RNS_PRIME_BITS'd785839955, `RNS_PRIME_BITS'd514404981, `RNS_PRIME_BITS'd1060123773, `RNS_PRIME_BITS'd1370482996, `RNS_PRIME_BITS'd1714034529, `RNS_PRIME_BITS'd176593021},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd1283744391, `RNS_PRIME_BITS'd392543978, `RNS_PRIME_BITS'd1911549448, `RNS_PRIME_BITS'd2142150955, `RNS_PRIME_BITS'd1226920252, `RNS_PRIME_BITS'd777751900, `RNS_PRIME_BITS'd624056478, `RNS_PRIME_BITS'd370579046, `RNS_PRIME_BITS'd204003667, `RNS_PRIME_BITS'd1425279212},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd863544926, `RNS_PRIME_BITS'd1129965629, `RNS_PRIME_BITS'd493869466, `RNS_PRIME_BITS'd2016533256, `RNS_PRIME_BITS'd2052423864, `RNS_PRIME_BITS'd128819871, `RNS_PRIME_BITS'd1269093335, `RNS_PRIME_BITS'd395823824, `RNS_PRIME_BITS'd1372360357, `RNS_PRIME_BITS'd432204286},
			'{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd1625556344, `RNS_PRIME_BITS'd403856286, `RNS_PRIME_BITS'd801996979, `RNS_PRIME_BITS'd1745818034, `RNS_PRIME_BITS'd1786207842, `RNS_PRIME_BITS'd736030319, `RNS_PRIME_BITS'd145225363, `RNS_PRIME_BITS'd275367179, `RNS_PRIME_BITS'd423711716, `RNS_PRIME_BITS'd802666385},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1105708626, `RNS_PRIME_BITS'd1726477570, `RNS_PRIME_BITS'd1574582621, `RNS_PRIME_BITS'd1199556620, `RNS_PRIME_BITS'd94276007, `RNS_PRIME_BITS'd1376820646, `RNS_PRIME_BITS'd17603037, `RNS_PRIME_BITS'd690382849, `RNS_PRIME_BITS'd2125518510, `RNS_PRIME_BITS'd305496598},
			'{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd1602274014, `RNS_PRIME_BITS'd1690084490, `RNS_PRIME_BITS'd1639860634, `RNS_PRIME_BITS'd1010974170, `RNS_PRIME_BITS'd661219551, `RNS_PRIME_BITS'd742474558, `RNS_PRIME_BITS'd1992932969, `RNS_PRIME_BITS'd1430056885, `RNS_PRIME_BITS'd227830247, `RNS_PRIME_BITS'd373164937},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1812739649, `RNS_PRIME_BITS'd1560593645, `RNS_PRIME_BITS'd228624354, `RNS_PRIME_BITS'd194524984, `RNS_PRIME_BITS'd252623462, `RNS_PRIME_BITS'd1008775490, `RNS_PRIME_BITS'd1973374751, `RNS_PRIME_BITS'd247231099, `RNS_PRIME_BITS'd989702289, `RNS_PRIME_BITS'd1998146343},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd726222268, `RNS_PRIME_BITS'd536389781, `RNS_PRIME_BITS'd1828738682, `RNS_PRIME_BITS'd1222472677, `RNS_PRIME_BITS'd1708734274, `RNS_PRIME_BITS'd1550286765, `RNS_PRIME_BITS'd1730816265, `RNS_PRIME_BITS'd508743819, `RNS_PRIME_BITS'd520970781, `RNS_PRIME_BITS'd1664611751},
			'{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd814240943, `RNS_PRIME_BITS'd66070744, `RNS_PRIME_BITS'd912999066, `RNS_PRIME_BITS'd1436211854, `RNS_PRIME_BITS'd1626275614, `RNS_PRIME_BITS'd303149686, `RNS_PRIME_BITS'd460768857, `RNS_PRIME_BITS'd1348884882, `RNS_PRIME_BITS'd1906010972, `RNS_PRIME_BITS'd556643362},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd742982649, `RNS_PRIME_BITS'd1425847407, `RNS_PRIME_BITS'd390431430, `RNS_PRIME_BITS'd1328059674, `RNS_PRIME_BITS'd570420539, `RNS_PRIME_BITS'd43469897, `RNS_PRIME_BITS'd1950964428, `RNS_PRIME_BITS'd643267493, `RNS_PRIME_BITS'd1108649918, `RNS_PRIME_BITS'd1008002272},
			'{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd996770076, `RNS_PRIME_BITS'd325882575, `RNS_PRIME_BITS'd1627184586, `RNS_PRIME_BITS'd205492666, `RNS_PRIME_BITS'd1643862925, `RNS_PRIME_BITS'd1793949804, `RNS_PRIME_BITS'd1920323117, `RNS_PRIME_BITS'd111054384, `RNS_PRIME_BITS'd1683505931, `RNS_PRIME_BITS'd1339474593},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd27672876, `RNS_PRIME_BITS'd1631145047, `RNS_PRIME_BITS'd1885928167, `RNS_PRIME_BITS'd629348003, `RNS_PRIME_BITS'd85973598, `RNS_PRIME_BITS'd2026186310, `RNS_PRIME_BITS'd335064443, `RNS_PRIME_BITS'd324888245, `RNS_PRIME_BITS'd1588230931, `RNS_PRIME_BITS'd313525161},
			'{`RNS_PRIME_BITS'd180, `RNS_PRIME_BITS'd290980759, `RNS_PRIME_BITS'd925640860, `RNS_PRIME_BITS'd1145801701, `RNS_PRIME_BITS'd1720573207, `RNS_PRIME_BITS'd1750329596, `RNS_PRIME_BITS'd785642955, `RNS_PRIME_BITS'd1887995987, `RNS_PRIME_BITS'd1625278573, `RNS_PRIME_BITS'd80813475, `RNS_PRIME_BITS'd953404240},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd1290020475, `RNS_PRIME_BITS'd1919566938, `RNS_PRIME_BITS'd2124724934, `RNS_PRIME_BITS'd1543702301, `RNS_PRIME_BITS'd245439945, `RNS_PRIME_BITS'd1875590086, `RNS_PRIME_BITS'd1421922164, `RNS_PRIME_BITS'd1979857703, `RNS_PRIME_BITS'd1094792709, `RNS_PRIME_BITS'd1556206507},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd333092724, `RNS_PRIME_BITS'd1951436064, `RNS_PRIME_BITS'd1135850590, `RNS_PRIME_BITS'd109454722, `RNS_PRIME_BITS'd216739934, `RNS_PRIME_BITS'd243989466, `RNS_PRIME_BITS'd1203261310, `RNS_PRIME_BITS'd758733881, `RNS_PRIME_BITS'd2070789561, `RNS_PRIME_BITS'd1696215523},
			'{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd1157123317, `RNS_PRIME_BITS'd1959724314, `RNS_PRIME_BITS'd948641442, `RNS_PRIME_BITS'd533660824, `RNS_PRIME_BITS'd1490620883, `RNS_PRIME_BITS'd540659115, `RNS_PRIME_BITS'd1017974019, `RNS_PRIME_BITS'd1724043246, `RNS_PRIME_BITS'd1719980946, `RNS_PRIME_BITS'd494425404},
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd15325996, `RNS_PRIME_BITS'd845742812, `RNS_PRIME_BITS'd996110387, `RNS_PRIME_BITS'd1333895523, `RNS_PRIME_BITS'd701744221, `RNS_PRIME_BITS'd1627895640, `RNS_PRIME_BITS'd1024699479, `RNS_PRIME_BITS'd1305064124, `RNS_PRIME_BITS'd1618567728, `RNS_PRIME_BITS'd1671651956},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd1302232967, `RNS_PRIME_BITS'd1518701377, `RNS_PRIME_BITS'd494721271, `RNS_PRIME_BITS'd496488456, `RNS_PRIME_BITS'd681852713, `RNS_PRIME_BITS'd1513193989, `RNS_PRIME_BITS'd1424915196, `RNS_PRIME_BITS'd1970475669, `RNS_PRIME_BITS'd1044199150, `RNS_PRIME_BITS'd1750380402},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd731603582, `RNS_PRIME_BITS'd1617525313, `RNS_PRIME_BITS'd856087701, `RNS_PRIME_BITS'd1707849750, `RNS_PRIME_BITS'd978340344, `RNS_PRIME_BITS'd425168302, `RNS_PRIME_BITS'd48108767, `RNS_PRIME_BITS'd412272618, `RNS_PRIME_BITS'd1067292332, `RNS_PRIME_BITS'd143175441},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd243159658, `RNS_PRIME_BITS'd1859710819, `RNS_PRIME_BITS'd279102314, `RNS_PRIME_BITS'd1736846096, `RNS_PRIME_BITS'd451617226, `RNS_PRIME_BITS'd176530023, `RNS_PRIME_BITS'd358278040, `RNS_PRIME_BITS'd556866622, `RNS_PRIME_BITS'd28708799, `RNS_PRIME_BITS'd4307079},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1217514340, `RNS_PRIME_BITS'd711842992, `RNS_PRIME_BITS'd498689010, `RNS_PRIME_BITS'd1261520405, `RNS_PRIME_BITS'd1728283132, `RNS_PRIME_BITS'd1197702349, `RNS_PRIME_BITS'd995124894, `RNS_PRIME_BITS'd1719909246, `RNS_PRIME_BITS'd2114687557, `RNS_PRIME_BITS'd1111271426},
			'{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd941726966, `RNS_PRIME_BITS'd4139816, `RNS_PRIME_BITS'd313983999, `RNS_PRIME_BITS'd1473489216, `RNS_PRIME_BITS'd1245157923, `RNS_PRIME_BITS'd290875422, `RNS_PRIME_BITS'd1826951809, `RNS_PRIME_BITS'd1310331238, `RNS_PRIME_BITS'd1841666462, `RNS_PRIME_BITS'd867524396},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd977138347, `RNS_PRIME_BITS'd1016520462, `RNS_PRIME_BITS'd1021398343, `RNS_PRIME_BITS'd619577642, `RNS_PRIME_BITS'd171881380, `RNS_PRIME_BITS'd1558258583, `RNS_PRIME_BITS'd780941068, `RNS_PRIME_BITS'd262755255, `RNS_PRIME_BITS'd2127218302, `RNS_PRIME_BITS'd691766545},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd124590189, `RNS_PRIME_BITS'd153024938, `RNS_PRIME_BITS'd380486293, `RNS_PRIME_BITS'd1625028206, `RNS_PRIME_BITS'd667652947, `RNS_PRIME_BITS'd1107446014, `RNS_PRIME_BITS'd1664507209, `RNS_PRIME_BITS'd950640035, `RNS_PRIME_BITS'd947949178, `RNS_PRIME_BITS'd1219988057},
			'{`RNS_PRIME_BITS'd54, `RNS_PRIME_BITS'd1476808599, `RNS_PRIME_BITS'd762239296, `RNS_PRIME_BITS'd1712403956, `RNS_PRIME_BITS'd657607857, `RNS_PRIME_BITS'd227939115, `RNS_PRIME_BITS'd1534771341, `RNS_PRIME_BITS'd141304030, `RNS_PRIME_BITS'd916948388, `RNS_PRIME_BITS'd1362103239, `RNS_PRIME_BITS'd1264765526},
			'{`RNS_PRIME_BITS'd69, `RNS_PRIME_BITS'd960556993, `RNS_PRIME_BITS'd2058637813, `RNS_PRIME_BITS'd1814282753, `RNS_PRIME_BITS'd862284988, `RNS_PRIME_BITS'd1687949847, `RNS_PRIME_BITS'd1116300621, `RNS_PRIME_BITS'd570004635, `RNS_PRIME_BITS'd1054747748, `RNS_PRIME_BITS'd1117355052, `RNS_PRIME_BITS'd922537397},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd2108497432, `RNS_PRIME_BITS'd299473228, `RNS_PRIME_BITS'd260764099, `RNS_PRIME_BITS'd49034613, `RNS_PRIME_BITS'd1771983436, `RNS_PRIME_BITS'd1591073326, `RNS_PRIME_BITS'd601369141, `RNS_PRIME_BITS'd168975701, `RNS_PRIME_BITS'd1886771897, `RNS_PRIME_BITS'd244786542},
			'{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd947536960, `RNS_PRIME_BITS'd1058553823, `RNS_PRIME_BITS'd494803513, `RNS_PRIME_BITS'd935961595, `RNS_PRIME_BITS'd1686724634, `RNS_PRIME_BITS'd1522670552, `RNS_PRIME_BITS'd1187826413, `RNS_PRIME_BITS'd587678567, `RNS_PRIME_BITS'd1912166830, `RNS_PRIME_BITS'd736574189},
			'{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd918251326, `RNS_PRIME_BITS'd1320750195, `RNS_PRIME_BITS'd2009641776, `RNS_PRIME_BITS'd331441599, `RNS_PRIME_BITS'd1017673839, `RNS_PRIME_BITS'd1212912172, `RNS_PRIME_BITS'd1922752404, `RNS_PRIME_BITS'd193404800, `RNS_PRIME_BITS'd1645799440, `RNS_PRIME_BITS'd1964889510},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd779152443, `RNS_PRIME_BITS'd1368543940, `RNS_PRIME_BITS'd1435061644, `RNS_PRIME_BITS'd229512241, `RNS_PRIME_BITS'd864840312, `RNS_PRIME_BITS'd2112701580, `RNS_PRIME_BITS'd1248112692, `RNS_PRIME_BITS'd10166037, `RNS_PRIME_BITS'd1380600983, `RNS_PRIME_BITS'd835715554},
			'{`RNS_PRIME_BITS'd238, `RNS_PRIME_BITS'd372364296, `RNS_PRIME_BITS'd1247659599, `RNS_PRIME_BITS'd1328891938, `RNS_PRIME_BITS'd2101541387, `RNS_PRIME_BITS'd720114338, `RNS_PRIME_BITS'd1815520558, `RNS_PRIME_BITS'd290109010, `RNS_PRIME_BITS'd12285042, `RNS_PRIME_BITS'd1346417431, `RNS_PRIME_BITS'd985589221},
			'{`RNS_PRIME_BITS'd32, `RNS_PRIME_BITS'd428316038, `RNS_PRIME_BITS'd1060816242, `RNS_PRIME_BITS'd862091863, `RNS_PRIME_BITS'd626573172, `RNS_PRIME_BITS'd1189997875, `RNS_PRIME_BITS'd450417019, `RNS_PRIME_BITS'd1734779829, `RNS_PRIME_BITS'd840243228, `RNS_PRIME_BITS'd166699489, `RNS_PRIME_BITS'd2143626148},
			'{`RNS_PRIME_BITS'd66, `RNS_PRIME_BITS'd1690699219, `RNS_PRIME_BITS'd1342201975, `RNS_PRIME_BITS'd415129330, `RNS_PRIME_BITS'd199965666, `RNS_PRIME_BITS'd396930850, `RNS_PRIME_BITS'd581327703, `RNS_PRIME_BITS'd414612647, `RNS_PRIME_BITS'd2083879465, `RNS_PRIME_BITS'd967877891, `RNS_PRIME_BITS'd134641468},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd2110307687, `RNS_PRIME_BITS'd450065239, `RNS_PRIME_BITS'd169957262, `RNS_PRIME_BITS'd318294795, `RNS_PRIME_BITS'd1382951105, `RNS_PRIME_BITS'd575570274, `RNS_PRIME_BITS'd1945860630, `RNS_PRIME_BITS'd1693211385, `RNS_PRIME_BITS'd1667450617, `RNS_PRIME_BITS'd955927744},
			'{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd1044891920, `RNS_PRIME_BITS'd1275633816, `RNS_PRIME_BITS'd1378358372, `RNS_PRIME_BITS'd1820699646, `RNS_PRIME_BITS'd1091440374, `RNS_PRIME_BITS'd2071157266, `RNS_PRIME_BITS'd1829417766, `RNS_PRIME_BITS'd89995327, `RNS_PRIME_BITS'd1725247476, `RNS_PRIME_BITS'd866796888},
			'{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd125990748, `RNS_PRIME_BITS'd499210037, `RNS_PRIME_BITS'd1055036707, `RNS_PRIME_BITS'd697936328, `RNS_PRIME_BITS'd1013996455, `RNS_PRIME_BITS'd591245625, `RNS_PRIME_BITS'd1187657455, `RNS_PRIME_BITS'd1898585489, `RNS_PRIME_BITS'd1050059250, `RNS_PRIME_BITS'd589451478},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd1762419996, `RNS_PRIME_BITS'd551707784, `RNS_PRIME_BITS'd1837146053, `RNS_PRIME_BITS'd789563477, `RNS_PRIME_BITS'd1762993140, `RNS_PRIME_BITS'd1797040315, `RNS_PRIME_BITS'd217372707, `RNS_PRIME_BITS'd374270343, `RNS_PRIME_BITS'd52129640, `RNS_PRIME_BITS'd295336306},
			'{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd253639859, `RNS_PRIME_BITS'd1076458040, `RNS_PRIME_BITS'd1128822673, `RNS_PRIME_BITS'd1483027350, `RNS_PRIME_BITS'd166126037, `RNS_PRIME_BITS'd662770625, `RNS_PRIME_BITS'd495773426, `RNS_PRIME_BITS'd2102707159, `RNS_PRIME_BITS'd296258777, `RNS_PRIME_BITS'd572957612},
			'{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd28576442, `RNS_PRIME_BITS'd1800392802, `RNS_PRIME_BITS'd1553903129, `RNS_PRIME_BITS'd1825458488, `RNS_PRIME_BITS'd1774013178, `RNS_PRIME_BITS'd813190193, `RNS_PRIME_BITS'd2127917048, `RNS_PRIME_BITS'd22041796, `RNS_PRIME_BITS'd1648387143, `RNS_PRIME_BITS'd1148697663},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd953850284, `RNS_PRIME_BITS'd140868616, `RNS_PRIME_BITS'd889981975, `RNS_PRIME_BITS'd1262581489, `RNS_PRIME_BITS'd1701391346, `RNS_PRIME_BITS'd883708958, `RNS_PRIME_BITS'd313585664, `RNS_PRIME_BITS'd1267682249, `RNS_PRIME_BITS'd1331216845, `RNS_PRIME_BITS'd927048052},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd355608994, `RNS_PRIME_BITS'd955780289, `RNS_PRIME_BITS'd269881985, `RNS_PRIME_BITS'd172876723, `RNS_PRIME_BITS'd1270243330, `RNS_PRIME_BITS'd613506468, `RNS_PRIME_BITS'd1891462904, `RNS_PRIME_BITS'd810512357, `RNS_PRIME_BITS'd554916618, `RNS_PRIME_BITS'd1103868672},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd571302931, `RNS_PRIME_BITS'd1058372862, `RNS_PRIME_BITS'd733508526, `RNS_PRIME_BITS'd967019763, `RNS_PRIME_BITS'd183441967, `RNS_PRIME_BITS'd976404709, `RNS_PRIME_BITS'd753601655, `RNS_PRIME_BITS'd1204654700, `RNS_PRIME_BITS'd1312266245, `RNS_PRIME_BITS'd241298613},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd775939505, `RNS_PRIME_BITS'd388499405, `RNS_PRIME_BITS'd924148638, `RNS_PRIME_BITS'd829105413, `RNS_PRIME_BITS'd1841635655, `RNS_PRIME_BITS'd959092768, `RNS_PRIME_BITS'd2043639771, `RNS_PRIME_BITS'd889685767, `RNS_PRIME_BITS'd160142765, `RNS_PRIME_BITS'd1465925103},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd2137835630, `RNS_PRIME_BITS'd1630642232, `RNS_PRIME_BITS'd1835327331, `RNS_PRIME_BITS'd303827008, `RNS_PRIME_BITS'd1937510308, `RNS_PRIME_BITS'd1001892870, `RNS_PRIME_BITS'd1184105923, `RNS_PRIME_BITS'd429394346, `RNS_PRIME_BITS'd1750753121, `RNS_PRIME_BITS'd1510096385},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd438668416, `RNS_PRIME_BITS'd442865527, `RNS_PRIME_BITS'd1773018651, `RNS_PRIME_BITS'd12789128, `RNS_PRIME_BITS'd1093820609, `RNS_PRIME_BITS'd1678966294, `RNS_PRIME_BITS'd52371623, `RNS_PRIME_BITS'd456791063, `RNS_PRIME_BITS'd801922940, `RNS_PRIME_BITS'd358501222},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd56929047, `RNS_PRIME_BITS'd1640141280, `RNS_PRIME_BITS'd68082040, `RNS_PRIME_BITS'd788328560, `RNS_PRIME_BITS'd653170079, `RNS_PRIME_BITS'd1538901594, `RNS_PRIME_BITS'd1820813304, `RNS_PRIME_BITS'd1541552150, `RNS_PRIME_BITS'd2076798616, `RNS_PRIME_BITS'd1441850245},
			'{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd1937725098, `RNS_PRIME_BITS'd1267001696, `RNS_PRIME_BITS'd733058130, `RNS_PRIME_BITS'd1553041679, `RNS_PRIME_BITS'd1634970318, `RNS_PRIME_BITS'd1541163766, `RNS_PRIME_BITS'd2013350457, `RNS_PRIME_BITS'd1694603161, `RNS_PRIME_BITS'd1227545592, `RNS_PRIME_BITS'd1402186930},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd831500109, `RNS_PRIME_BITS'd902929161, `RNS_PRIME_BITS'd1291235238, `RNS_PRIME_BITS'd1424507932, `RNS_PRIME_BITS'd476913892, `RNS_PRIME_BITS'd551316114, `RNS_PRIME_BITS'd476637886, `RNS_PRIME_BITS'd874386955, `RNS_PRIME_BITS'd1862806601, `RNS_PRIME_BITS'd1577901434},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1931392889, `RNS_PRIME_BITS'd1974498828, `RNS_PRIME_BITS'd450850943, `RNS_PRIME_BITS'd835327743, `RNS_PRIME_BITS'd125057386, `RNS_PRIME_BITS'd669245744, `RNS_PRIME_BITS'd1080019999, `RNS_PRIME_BITS'd611814508, `RNS_PRIME_BITS'd1731351620, `RNS_PRIME_BITS'd76983612},
			'{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd152049574, `RNS_PRIME_BITS'd2023773705, `RNS_PRIME_BITS'd110962637, `RNS_PRIME_BITS'd663796804, `RNS_PRIME_BITS'd1783124859, `RNS_PRIME_BITS'd1694610459, `RNS_PRIME_BITS'd1575031362, `RNS_PRIME_BITS'd1390089269, `RNS_PRIME_BITS'd1799987617, `RNS_PRIME_BITS'd489685295},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd1785890277, `RNS_PRIME_BITS'd739416543, `RNS_PRIME_BITS'd1059186330, `RNS_PRIME_BITS'd341091810, `RNS_PRIME_BITS'd1484422994, `RNS_PRIME_BITS'd962270263, `RNS_PRIME_BITS'd528875623, `RNS_PRIME_BITS'd1395267808, `RNS_PRIME_BITS'd731815571, `RNS_PRIME_BITS'd1282564241},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd298204622, `RNS_PRIME_BITS'd1821128942, `RNS_PRIME_BITS'd1123923466, `RNS_PRIME_BITS'd597296355, `RNS_PRIME_BITS'd284692885, `RNS_PRIME_BITS'd25333225, `RNS_PRIME_BITS'd1202166285, `RNS_PRIME_BITS'd1856015609, `RNS_PRIME_BITS'd1802548151, `RNS_PRIME_BITS'd1352876417},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd299794594, `RNS_PRIME_BITS'd1500094201, `RNS_PRIME_BITS'd1029270485, `RNS_PRIME_BITS'd1957189005, `RNS_PRIME_BITS'd1074382340, `RNS_PRIME_BITS'd682031018, `RNS_PRIME_BITS'd118828473, `RNS_PRIME_BITS'd540216927, `RNS_PRIME_BITS'd1702305861, `RNS_PRIME_BITS'd278042139},
			'{`RNS_PRIME_BITS'd86, `RNS_PRIME_BITS'd1540340409, `RNS_PRIME_BITS'd1062372187, `RNS_PRIME_BITS'd1128409765, `RNS_PRIME_BITS'd348779406, `RNS_PRIME_BITS'd1093591790, `RNS_PRIME_BITS'd1695755043, `RNS_PRIME_BITS'd1219055793, `RNS_PRIME_BITS'd1934040631, `RNS_PRIME_BITS'd1148397770, `RNS_PRIME_BITS'd291330641},
			'{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd1969032376, `RNS_PRIME_BITS'd1591717252, `RNS_PRIME_BITS'd1152159931, `RNS_PRIME_BITS'd2145300746, `RNS_PRIME_BITS'd848800218, `RNS_PRIME_BITS'd155936820, `RNS_PRIME_BITS'd1309965203, `RNS_PRIME_BITS'd121669610, `RNS_PRIME_BITS'd1496733764, `RNS_PRIME_BITS'd925031395},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd1504712853, `RNS_PRIME_BITS'd2114512934, `RNS_PRIME_BITS'd1855683509, `RNS_PRIME_BITS'd756444084, `RNS_PRIME_BITS'd804844185, `RNS_PRIME_BITS'd758136197, `RNS_PRIME_BITS'd511032546, `RNS_PRIME_BITS'd1614555499, `RNS_PRIME_BITS'd150822317, `RNS_PRIME_BITS'd1270100314},
			'{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd562924617, `RNS_PRIME_BITS'd1433534961, `RNS_PRIME_BITS'd257262409, `RNS_PRIME_BITS'd1236112613, `RNS_PRIME_BITS'd1584702211, `RNS_PRIME_BITS'd163863614, `RNS_PRIME_BITS'd1433891858, `RNS_PRIME_BITS'd1436025740, `RNS_PRIME_BITS'd513755285, `RNS_PRIME_BITS'd1865153309},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1745932387, `RNS_PRIME_BITS'd370990367, `RNS_PRIME_BITS'd1922181368, `RNS_PRIME_BITS'd1004335570, `RNS_PRIME_BITS'd906538739, `RNS_PRIME_BITS'd1725596490, `RNS_PRIME_BITS'd832071432, `RNS_PRIME_BITS'd1784145682, `RNS_PRIME_BITS'd2057455634, `RNS_PRIME_BITS'd1097306852},
			'{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd1773019225, `RNS_PRIME_BITS'd1229377751, `RNS_PRIME_BITS'd450722484, `RNS_PRIME_BITS'd508434771, `RNS_PRIME_BITS'd1803880500, `RNS_PRIME_BITS'd2127566149, `RNS_PRIME_BITS'd561799542, `RNS_PRIME_BITS'd287961602, `RNS_PRIME_BITS'd1631705977, `RNS_PRIME_BITS'd109580911}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd1603204325, `RNS_PRIME_BITS'd65919473, `RNS_PRIME_BITS'd274808067, `RNS_PRIME_BITS'd1837766162, `RNS_PRIME_BITS'd740791666, `RNS_PRIME_BITS'd1640991241, `RNS_PRIME_BITS'd1687453662, `RNS_PRIME_BITS'd8323732, `RNS_PRIME_BITS'd591156347, `RNS_PRIME_BITS'd1264580105},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd186173184, `RNS_PRIME_BITS'd1361649095, `RNS_PRIME_BITS'd216316379, `RNS_PRIME_BITS'd1435086423, `RNS_PRIME_BITS'd913383032, `RNS_PRIME_BITS'd2113961977, `RNS_PRIME_BITS'd1009888390, `RNS_PRIME_BITS'd1689229263, `RNS_PRIME_BITS'd1591570223, `RNS_PRIME_BITS'd1847755074},
			'{`RNS_PRIME_BITS'd202, `RNS_PRIME_BITS'd12257270, `RNS_PRIME_BITS'd1695801865, `RNS_PRIME_BITS'd924964826, `RNS_PRIME_BITS'd919037594, `RNS_PRIME_BITS'd1158448048, `RNS_PRIME_BITS'd1615395084, `RNS_PRIME_BITS'd599564329, `RNS_PRIME_BITS'd1527434235, `RNS_PRIME_BITS'd807879414, `RNS_PRIME_BITS'd1464521084},
			'{`RNS_PRIME_BITS'd179, `RNS_PRIME_BITS'd247723499, `RNS_PRIME_BITS'd1218950578, `RNS_PRIME_BITS'd1325661954, `RNS_PRIME_BITS'd1982623594, `RNS_PRIME_BITS'd12617824, `RNS_PRIME_BITS'd1412720003, `RNS_PRIME_BITS'd835315677, `RNS_PRIME_BITS'd136313712, `RNS_PRIME_BITS'd1468499845, `RNS_PRIME_BITS'd1158897717},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd450848040, `RNS_PRIME_BITS'd592100019, `RNS_PRIME_BITS'd89411169, `RNS_PRIME_BITS'd1593549479, `RNS_PRIME_BITS'd1292088992, `RNS_PRIME_BITS'd1454046901, `RNS_PRIME_BITS'd527549415, `RNS_PRIME_BITS'd1270195724, `RNS_PRIME_BITS'd711587904, `RNS_PRIME_BITS'd742393955},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1291797997, `RNS_PRIME_BITS'd1270275017, `RNS_PRIME_BITS'd1165101958, `RNS_PRIME_BITS'd1293961455, `RNS_PRIME_BITS'd229837467, `RNS_PRIME_BITS'd88844973, `RNS_PRIME_BITS'd926301664, `RNS_PRIME_BITS'd714062608, `RNS_PRIME_BITS'd2076359092, `RNS_PRIME_BITS'd213394685},
			'{`RNS_PRIME_BITS'd20, `RNS_PRIME_BITS'd1169895117, `RNS_PRIME_BITS'd669930362, `RNS_PRIME_BITS'd5807910, `RNS_PRIME_BITS'd822430567, `RNS_PRIME_BITS'd2044073075, `RNS_PRIME_BITS'd1683706468, `RNS_PRIME_BITS'd812387325, `RNS_PRIME_BITS'd1631486604, `RNS_PRIME_BITS'd1865632943, `RNS_PRIME_BITS'd2025513155},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1797775022, `RNS_PRIME_BITS'd1308276368, `RNS_PRIME_BITS'd332757079, `RNS_PRIME_BITS'd239199367, `RNS_PRIME_BITS'd372704973, `RNS_PRIME_BITS'd1007840873, `RNS_PRIME_BITS'd1398574369, `RNS_PRIME_BITS'd1661833533, `RNS_PRIME_BITS'd1314760340, `RNS_PRIME_BITS'd2075416387},
			'{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd2018737179, `RNS_PRIME_BITS'd177362100, `RNS_PRIME_BITS'd1243823238, `RNS_PRIME_BITS'd1522000526, `RNS_PRIME_BITS'd314610333, `RNS_PRIME_BITS'd789740479, `RNS_PRIME_BITS'd1400047360, `RNS_PRIME_BITS'd502884766, `RNS_PRIME_BITS'd1553035696, `RNS_PRIME_BITS'd651536648},
			'{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd552444074, `RNS_PRIME_BITS'd1500389490, `RNS_PRIME_BITS'd1012168146, `RNS_PRIME_BITS'd1026954809, `RNS_PRIME_BITS'd2123068850, `RNS_PRIME_BITS'd161104410, `RNS_PRIME_BITS'd1463382507, `RNS_PRIME_BITS'd928257670, `RNS_PRIME_BITS'd832574682, `RNS_PRIME_BITS'd411868450},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd639946122, `RNS_PRIME_BITS'd1341759485, `RNS_PRIME_BITS'd1378190757, `RNS_PRIME_BITS'd1341919726, `RNS_PRIME_BITS'd1538049989, `RNS_PRIME_BITS'd459002246, `RNS_PRIME_BITS'd772327900, `RNS_PRIME_BITS'd493083855, `RNS_PRIME_BITS'd811041990, `RNS_PRIME_BITS'd1336643866},
			'{`RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd2126183905, `RNS_PRIME_BITS'd188678037, `RNS_PRIME_BITS'd805777536, `RNS_PRIME_BITS'd1743013868, `RNS_PRIME_BITS'd1084291413, `RNS_PRIME_BITS'd1712703081, `RNS_PRIME_BITS'd25420016, `RNS_PRIME_BITS'd2066467423, `RNS_PRIME_BITS'd305033547, `RNS_PRIME_BITS'd610674220},
			'{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd152066605, `RNS_PRIME_BITS'd636894190, `RNS_PRIME_BITS'd1943582733, `RNS_PRIME_BITS'd1070421290, `RNS_PRIME_BITS'd2095770421, `RNS_PRIME_BITS'd1105205300, `RNS_PRIME_BITS'd880862598, `RNS_PRIME_BITS'd1864718971, `RNS_PRIME_BITS'd808865573, `RNS_PRIME_BITS'd1803539214},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd1273359706, `RNS_PRIME_BITS'd68162432, `RNS_PRIME_BITS'd22716372, `RNS_PRIME_BITS'd1405249091, `RNS_PRIME_BITS'd1506397445, `RNS_PRIME_BITS'd486885848, `RNS_PRIME_BITS'd500596407, `RNS_PRIME_BITS'd632812140, `RNS_PRIME_BITS'd1598457887, `RNS_PRIME_BITS'd313681499},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd350062283, `RNS_PRIME_BITS'd17496022, `RNS_PRIME_BITS'd1596533811, `RNS_PRIME_BITS'd446315255, `RNS_PRIME_BITS'd1431248847, `RNS_PRIME_BITS'd906992474, `RNS_PRIME_BITS'd453321261, `RNS_PRIME_BITS'd1554627360, `RNS_PRIME_BITS'd77942201, `RNS_PRIME_BITS'd2002489505},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd2127302935, `RNS_PRIME_BITS'd2042009268, `RNS_PRIME_BITS'd352985053, `RNS_PRIME_BITS'd303002740, `RNS_PRIME_BITS'd2001007184, `RNS_PRIME_BITS'd641353728, `RNS_PRIME_BITS'd135918769, `RNS_PRIME_BITS'd439702740, `RNS_PRIME_BITS'd880721004, `RNS_PRIME_BITS'd1311622039},
			'{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd846272909, `RNS_PRIME_BITS'd1393384121, `RNS_PRIME_BITS'd2005559565, `RNS_PRIME_BITS'd1015410496, `RNS_PRIME_BITS'd1621639016, `RNS_PRIME_BITS'd963656143, `RNS_PRIME_BITS'd647787250, `RNS_PRIME_BITS'd504170809, `RNS_PRIME_BITS'd108035381, `RNS_PRIME_BITS'd501262205},
			'{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd1723349031, `RNS_PRIME_BITS'd688117755, `RNS_PRIME_BITS'd969735708, `RNS_PRIME_BITS'd1270498877, `RNS_PRIME_BITS'd57863878, `RNS_PRIME_BITS'd1877837595, `RNS_PRIME_BITS'd1627361466, `RNS_PRIME_BITS'd1784089160, `RNS_PRIME_BITS'd1616617931, `RNS_PRIME_BITS'd972067593},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd272417344, `RNS_PRIME_BITS'd1676768779, `RNS_PRIME_BITS'd737764576, `RNS_PRIME_BITS'd244397223, `RNS_PRIME_BITS'd1843251163, `RNS_PRIME_BITS'd1578410639, `RNS_PRIME_BITS'd316057477, `RNS_PRIME_BITS'd74084405, `RNS_PRIME_BITS'd412585241, `RNS_PRIME_BITS'd992453593},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd622014856, `RNS_PRIME_BITS'd673632700, `RNS_PRIME_BITS'd1553140577, `RNS_PRIME_BITS'd1473701546, `RNS_PRIME_BITS'd669889421, `RNS_PRIME_BITS'd43212541, `RNS_PRIME_BITS'd393392585, `RNS_PRIME_BITS'd1248030717, `RNS_PRIME_BITS'd1483349072, `RNS_PRIME_BITS'd2012470289},
			'{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd1815539687, `RNS_PRIME_BITS'd265765934, `RNS_PRIME_BITS'd954158022, `RNS_PRIME_BITS'd1454637123, `RNS_PRIME_BITS'd1888433019, `RNS_PRIME_BITS'd556442916, `RNS_PRIME_BITS'd553695888, `RNS_PRIME_BITS'd731363658, `RNS_PRIME_BITS'd210890704, `RNS_PRIME_BITS'd448889365},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd1513104184, `RNS_PRIME_BITS'd1453656356, `RNS_PRIME_BITS'd352694716, `RNS_PRIME_BITS'd2124947579, `RNS_PRIME_BITS'd484859594, `RNS_PRIME_BITS'd1904817924, `RNS_PRIME_BITS'd531797433, `RNS_PRIME_BITS'd962191838, `RNS_PRIME_BITS'd173514477, `RNS_PRIME_BITS'd1081286762},
			'{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd1734848078, `RNS_PRIME_BITS'd1742126284, `RNS_PRIME_BITS'd1612799781, `RNS_PRIME_BITS'd1564126038, `RNS_PRIME_BITS'd1132105068, `RNS_PRIME_BITS'd1957714917, `RNS_PRIME_BITS'd1741188534, `RNS_PRIME_BITS'd2012981777, `RNS_PRIME_BITS'd1272574458, `RNS_PRIME_BITS'd1022674347},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd1713016986, `RNS_PRIME_BITS'd712034409, `RNS_PRIME_BITS'd1342535935, `RNS_PRIME_BITS'd806010628, `RNS_PRIME_BITS'd963904170, `RNS_PRIME_BITS'd2101710850, `RNS_PRIME_BITS'd1654720077, `RNS_PRIME_BITS'd1853015878, `RNS_PRIME_BITS'd847821514, `RNS_PRIME_BITS'd173312846},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1807451681, `RNS_PRIME_BITS'd766838182, `RNS_PRIME_BITS'd1820672985, `RNS_PRIME_BITS'd355794089, `RNS_PRIME_BITS'd537553304, `RNS_PRIME_BITS'd1486416655, `RNS_PRIME_BITS'd1218013184, `RNS_PRIME_BITS'd1403447957, `RNS_PRIME_BITS'd302458652, `RNS_PRIME_BITS'd1554874283},
			'{`RNS_PRIME_BITS'd201, `RNS_PRIME_BITS'd606675239, `RNS_PRIME_BITS'd655824039, `RNS_PRIME_BITS'd874995568, `RNS_PRIME_BITS'd952326726, `RNS_PRIME_BITS'd1629549131, `RNS_PRIME_BITS'd678219044, `RNS_PRIME_BITS'd581116066, `RNS_PRIME_BITS'd909148296, `RNS_PRIME_BITS'd354715650, `RNS_PRIME_BITS'd1498775119},
			'{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd2039986956, `RNS_PRIME_BITS'd189066492, `RNS_PRIME_BITS'd727879070, `RNS_PRIME_BITS'd1984847273, `RNS_PRIME_BITS'd1608976089, `RNS_PRIME_BITS'd952654308, `RNS_PRIME_BITS'd1919565238, `RNS_PRIME_BITS'd1768747349, `RNS_PRIME_BITS'd1553704756, `RNS_PRIME_BITS'd1286675246},
			'{`RNS_PRIME_BITS'd160, `RNS_PRIME_BITS'd1088284398, `RNS_PRIME_BITS'd455656220, `RNS_PRIME_BITS'd253795628, `RNS_PRIME_BITS'd324532434, `RNS_PRIME_BITS'd1915378432, `RNS_PRIME_BITS'd657441659, `RNS_PRIME_BITS'd733450532, `RNS_PRIME_BITS'd1553149242, `RNS_PRIME_BITS'd103240049, `RNS_PRIME_BITS'd427886149},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd473098862, `RNS_PRIME_BITS'd137263828, `RNS_PRIME_BITS'd781856744, `RNS_PRIME_BITS'd1071571904, `RNS_PRIME_BITS'd883343976, `RNS_PRIME_BITS'd1922990766, `RNS_PRIME_BITS'd763483046, `RNS_PRIME_BITS'd240132974, `RNS_PRIME_BITS'd988363126, `RNS_PRIME_BITS'd190822907},
			'{`RNS_PRIME_BITS'd51, `RNS_PRIME_BITS'd914465651, `RNS_PRIME_BITS'd2058657397, `RNS_PRIME_BITS'd805880414, `RNS_PRIME_BITS'd136739468, `RNS_PRIME_BITS'd161493818, `RNS_PRIME_BITS'd268222657, `RNS_PRIME_BITS'd744942199, `RNS_PRIME_BITS'd1006473070, `RNS_PRIME_BITS'd1792394963, `RNS_PRIME_BITS'd232360598},
			'{`RNS_PRIME_BITS'd201, `RNS_PRIME_BITS'd2096115588, `RNS_PRIME_BITS'd904472948, `RNS_PRIME_BITS'd718360342, `RNS_PRIME_BITS'd403143559, `RNS_PRIME_BITS'd623099712, `RNS_PRIME_BITS'd2028461057, `RNS_PRIME_BITS'd1164870067, `RNS_PRIME_BITS'd1171189660, `RNS_PRIME_BITS'd501246767, `RNS_PRIME_BITS'd362547244},
			'{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd1322540935, `RNS_PRIME_BITS'd991977741, `RNS_PRIME_BITS'd862256936, `RNS_PRIME_BITS'd1793759105, `RNS_PRIME_BITS'd2048984760, `RNS_PRIME_BITS'd844727131, `RNS_PRIME_BITS'd235637592, `RNS_PRIME_BITS'd1804095556, `RNS_PRIME_BITS'd1941061966, `RNS_PRIME_BITS'd730684490},
			'{`RNS_PRIME_BITS'd204, `RNS_PRIME_BITS'd1731970645, `RNS_PRIME_BITS'd376926700, `RNS_PRIME_BITS'd1324443849, `RNS_PRIME_BITS'd808349914, `RNS_PRIME_BITS'd1613759621, `RNS_PRIME_BITS'd1884571882, `RNS_PRIME_BITS'd1625034437, `RNS_PRIME_BITS'd1848691393, `RNS_PRIME_BITS'd1962644574, `RNS_PRIME_BITS'd111810179},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd982313297, `RNS_PRIME_BITS'd1528940813, `RNS_PRIME_BITS'd1719388342, `RNS_PRIME_BITS'd1835202582, `RNS_PRIME_BITS'd1124799224, `RNS_PRIME_BITS'd1884080980, `RNS_PRIME_BITS'd1100309796, `RNS_PRIME_BITS'd1373114842, `RNS_PRIME_BITS'd344450970, `RNS_PRIME_BITS'd1061905760},
			'{`RNS_PRIME_BITS'd37, `RNS_PRIME_BITS'd113206552, `RNS_PRIME_BITS'd504986617, `RNS_PRIME_BITS'd371023110, `RNS_PRIME_BITS'd898553402, `RNS_PRIME_BITS'd575585562, `RNS_PRIME_BITS'd971339727, `RNS_PRIME_BITS'd824720065, `RNS_PRIME_BITS'd1688894077, `RNS_PRIME_BITS'd738346276, `RNS_PRIME_BITS'd1826479659},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd111878755, `RNS_PRIME_BITS'd1753175843, `RNS_PRIME_BITS'd1644568585, `RNS_PRIME_BITS'd1875922142, `RNS_PRIME_BITS'd1916309420, `RNS_PRIME_BITS'd1621347938, `RNS_PRIME_BITS'd1139633610, `RNS_PRIME_BITS'd1744338679, `RNS_PRIME_BITS'd1677534120, `RNS_PRIME_BITS'd521646467},
			'{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd610334054, `RNS_PRIME_BITS'd522703511, `RNS_PRIME_BITS'd844107222, `RNS_PRIME_BITS'd1170307646, `RNS_PRIME_BITS'd781087817, `RNS_PRIME_BITS'd818749035, `RNS_PRIME_BITS'd1638328007, `RNS_PRIME_BITS'd139534469, `RNS_PRIME_BITS'd1675670457, `RNS_PRIME_BITS'd474019076},
			'{`RNS_PRIME_BITS'd220, `RNS_PRIME_BITS'd541943610, `RNS_PRIME_BITS'd1311369917, `RNS_PRIME_BITS'd1908830868, `RNS_PRIME_BITS'd1300698844, `RNS_PRIME_BITS'd792043968, `RNS_PRIME_BITS'd1074677154, `RNS_PRIME_BITS'd947447869, `RNS_PRIME_BITS'd1666011340, `RNS_PRIME_BITS'd1463249565, `RNS_PRIME_BITS'd1119252872},
			'{`RNS_PRIME_BITS'd108, `RNS_PRIME_BITS'd956039615, `RNS_PRIME_BITS'd956381469, `RNS_PRIME_BITS'd583861817, `RNS_PRIME_BITS'd216531863, `RNS_PRIME_BITS'd1936573648, `RNS_PRIME_BITS'd2082974379, `RNS_PRIME_BITS'd2043905695, `RNS_PRIME_BITS'd1677884562, `RNS_PRIME_BITS'd992290593, `RNS_PRIME_BITS'd1529743842},
			'{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd1477803090, `RNS_PRIME_BITS'd1032297940, `RNS_PRIME_BITS'd1586157794, `RNS_PRIME_BITS'd1150504407, `RNS_PRIME_BITS'd765191635, `RNS_PRIME_BITS'd1936347998, `RNS_PRIME_BITS'd1490488316, `RNS_PRIME_BITS'd1175454414, `RNS_PRIME_BITS'd93829243, `RNS_PRIME_BITS'd1896501211},
			'{`RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd461269078, `RNS_PRIME_BITS'd201113189, `RNS_PRIME_BITS'd878151991, `RNS_PRIME_BITS'd1445947677, `RNS_PRIME_BITS'd1124795371, `RNS_PRIME_BITS'd818361039, `RNS_PRIME_BITS'd616303522, `RNS_PRIME_BITS'd1351968718, `RNS_PRIME_BITS'd1688730493, `RNS_PRIME_BITS'd2138880510},
			'{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd1208753729, `RNS_PRIME_BITS'd1986355259, `RNS_PRIME_BITS'd1353056259, `RNS_PRIME_BITS'd1719362313, `RNS_PRIME_BITS'd1970998302, `RNS_PRIME_BITS'd645272983, `RNS_PRIME_BITS'd978038662, `RNS_PRIME_BITS'd218337555, `RNS_PRIME_BITS'd1354571538, `RNS_PRIME_BITS'd713290017},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1017201423, `RNS_PRIME_BITS'd1619158017, `RNS_PRIME_BITS'd242875336, `RNS_PRIME_BITS'd403404819, `RNS_PRIME_BITS'd1400472835, `RNS_PRIME_BITS'd1756305608, `RNS_PRIME_BITS'd224881107, `RNS_PRIME_BITS'd1822798509, `RNS_PRIME_BITS'd961773138, `RNS_PRIME_BITS'd42454799},
			'{`RNS_PRIME_BITS'd127, `RNS_PRIME_BITS'd1737297970, `RNS_PRIME_BITS'd984441342, `RNS_PRIME_BITS'd978434081, `RNS_PRIME_BITS'd847499455, `RNS_PRIME_BITS'd263583318, `RNS_PRIME_BITS'd74992572, `RNS_PRIME_BITS'd1405678032, `RNS_PRIME_BITS'd1634657955, `RNS_PRIME_BITS'd1970857258, `RNS_PRIME_BITS'd981970991},
			'{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd2115091484, `RNS_PRIME_BITS'd165819299, `RNS_PRIME_BITS'd1419452784, `RNS_PRIME_BITS'd1955111196, `RNS_PRIME_BITS'd887497656, `RNS_PRIME_BITS'd305924393, `RNS_PRIME_BITS'd681954192, `RNS_PRIME_BITS'd1197700756, `RNS_PRIME_BITS'd264847438, `RNS_PRIME_BITS'd655490932},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd1732824386, `RNS_PRIME_BITS'd1142918605, `RNS_PRIME_BITS'd998801000, `RNS_PRIME_BITS'd1065530836, `RNS_PRIME_BITS'd237589369, `RNS_PRIME_BITS'd1620756877, `RNS_PRIME_BITS'd1878216831, `RNS_PRIME_BITS'd175422217, `RNS_PRIME_BITS'd1183132296, `RNS_PRIME_BITS'd1254449368},
			'{`RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd1081714830, `RNS_PRIME_BITS'd1980070825, `RNS_PRIME_BITS'd474673979, `RNS_PRIME_BITS'd313529963, `RNS_PRIME_BITS'd1827918201, `RNS_PRIME_BITS'd921018151, `RNS_PRIME_BITS'd1521233270, `RNS_PRIME_BITS'd1351762336, `RNS_PRIME_BITS'd149885184, `RNS_PRIME_BITS'd1618129381},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd338532842, `RNS_PRIME_BITS'd996511467, `RNS_PRIME_BITS'd1414400546, `RNS_PRIME_BITS'd2033404364, `RNS_PRIME_BITS'd2085804256, `RNS_PRIME_BITS'd1384162913, `RNS_PRIME_BITS'd1283083405, `RNS_PRIME_BITS'd2101513577, `RNS_PRIME_BITS'd96291307, `RNS_PRIME_BITS'd1627900336},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1504005917, `RNS_PRIME_BITS'd1486252548, `RNS_PRIME_BITS'd1371345878, `RNS_PRIME_BITS'd1200364540, `RNS_PRIME_BITS'd1287231700, `RNS_PRIME_BITS'd685020834, `RNS_PRIME_BITS'd405022461, `RNS_PRIME_BITS'd287768292, `RNS_PRIME_BITS'd1407969603, `RNS_PRIME_BITS'd2034627102},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd336451252, `RNS_PRIME_BITS'd110663629, `RNS_PRIME_BITS'd1740542532, `RNS_PRIME_BITS'd1994911148, `RNS_PRIME_BITS'd1863416939, `RNS_PRIME_BITS'd1280488260, `RNS_PRIME_BITS'd1701572421, `RNS_PRIME_BITS'd234743337, `RNS_PRIME_BITS'd1364767155, `RNS_PRIME_BITS'd1891494426},
			'{`RNS_PRIME_BITS'd22, `RNS_PRIME_BITS'd1776383843, `RNS_PRIME_BITS'd1158149199, `RNS_PRIME_BITS'd2017935920, `RNS_PRIME_BITS'd681467210, `RNS_PRIME_BITS'd780449965, `RNS_PRIME_BITS'd1422874265, `RNS_PRIME_BITS'd1218656160, `RNS_PRIME_BITS'd1478054451, `RNS_PRIME_BITS'd1682385595, `RNS_PRIME_BITS'd1209578678},
			'{`RNS_PRIME_BITS'd224, `RNS_PRIME_BITS'd2077006510, `RNS_PRIME_BITS'd695292991, `RNS_PRIME_BITS'd1059719590, `RNS_PRIME_BITS'd605266679, `RNS_PRIME_BITS'd299525225, `RNS_PRIME_BITS'd1717312729, `RNS_PRIME_BITS'd1543238019, `RNS_PRIME_BITS'd1436542827, `RNS_PRIME_BITS'd354162670, `RNS_PRIME_BITS'd454228504},
			'{`RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd777548303, `RNS_PRIME_BITS'd1767566955, `RNS_PRIME_BITS'd1284399228, `RNS_PRIME_BITS'd374133047, `RNS_PRIME_BITS'd1728345861, `RNS_PRIME_BITS'd1723195018, `RNS_PRIME_BITS'd1884046438, `RNS_PRIME_BITS'd1754481078, `RNS_PRIME_BITS'd78176546, `RNS_PRIME_BITS'd1405885564},
			'{`RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd1218483088, `RNS_PRIME_BITS'd74197350, `RNS_PRIME_BITS'd1917577004, `RNS_PRIME_BITS'd853540546, `RNS_PRIME_BITS'd1687383187, `RNS_PRIME_BITS'd2121330918, `RNS_PRIME_BITS'd1464955074, `RNS_PRIME_BITS'd759111785, `RNS_PRIME_BITS'd499644838, `RNS_PRIME_BITS'd710056053},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd1627798984, `RNS_PRIME_BITS'd925489499, `RNS_PRIME_BITS'd1623026685, `RNS_PRIME_BITS'd1938368762, `RNS_PRIME_BITS'd847070973, `RNS_PRIME_BITS'd1009799294, `RNS_PRIME_BITS'd1092668911, `RNS_PRIME_BITS'd19471505, `RNS_PRIME_BITS'd1839466173, `RNS_PRIME_BITS'd943919978},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1651987507, `RNS_PRIME_BITS'd308249625, `RNS_PRIME_BITS'd1147499924, `RNS_PRIME_BITS'd2046226877, `RNS_PRIME_BITS'd1700950713, `RNS_PRIME_BITS'd158968243, `RNS_PRIME_BITS'd1079213256, `RNS_PRIME_BITS'd1210942849, `RNS_PRIME_BITS'd1044104614, `RNS_PRIME_BITS'd1523849772},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd1433571549, `RNS_PRIME_BITS'd1566402292, `RNS_PRIME_BITS'd1841937957, `RNS_PRIME_BITS'd841374354, `RNS_PRIME_BITS'd51962549, `RNS_PRIME_BITS'd365026728, `RNS_PRIME_BITS'd17465727, `RNS_PRIME_BITS'd156906670, `RNS_PRIME_BITS'd1326637496, `RNS_PRIME_BITS'd670102719},
			'{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd1413979918, `RNS_PRIME_BITS'd188594269, `RNS_PRIME_BITS'd1831665972, `RNS_PRIME_BITS'd435747488, `RNS_PRIME_BITS'd1819450262, `RNS_PRIME_BITS'd1997875700, `RNS_PRIME_BITS'd777068210, `RNS_PRIME_BITS'd1202969192, `RNS_PRIME_BITS'd1362298696, `RNS_PRIME_BITS'd1263722878},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd551534351, `RNS_PRIME_BITS'd1896452170, `RNS_PRIME_BITS'd14636061, `RNS_PRIME_BITS'd1125495787, `RNS_PRIME_BITS'd2054139093, `RNS_PRIME_BITS'd1271566322, `RNS_PRIME_BITS'd1772482830, `RNS_PRIME_BITS'd1067690016, `RNS_PRIME_BITS'd865825036, `RNS_PRIME_BITS'd2050728258},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd1020882969, `RNS_PRIME_BITS'd858740119, `RNS_PRIME_BITS'd1040641671, `RNS_PRIME_BITS'd881138829, `RNS_PRIME_BITS'd297846696, `RNS_PRIME_BITS'd1921235899, `RNS_PRIME_BITS'd1496358970, `RNS_PRIME_BITS'd2123900040, `RNS_PRIME_BITS'd83607084, `RNS_PRIME_BITS'd156242963},
			'{`RNS_PRIME_BITS'd254, `RNS_PRIME_BITS'd1631323419, `RNS_PRIME_BITS'd1257032888, `RNS_PRIME_BITS'd1319197367, `RNS_PRIME_BITS'd1017172497, `RNS_PRIME_BITS'd1654427493, `RNS_PRIME_BITS'd1187235285, `RNS_PRIME_BITS'd1763683085, `RNS_PRIME_BITS'd1351866670, `RNS_PRIME_BITS'd5543773, `RNS_PRIME_BITS'd517243402},
			'{`RNS_PRIME_BITS'd167, `RNS_PRIME_BITS'd594869135, `RNS_PRIME_BITS'd1093422681, `RNS_PRIME_BITS'd1252710418, `RNS_PRIME_BITS'd1946306598, `RNS_PRIME_BITS'd292446400, `RNS_PRIME_BITS'd452576692, `RNS_PRIME_BITS'd1017142583, `RNS_PRIME_BITS'd490307155, `RNS_PRIME_BITS'd2003962294, `RNS_PRIME_BITS'd737954074},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1851847551, `RNS_PRIME_BITS'd1330922623, `RNS_PRIME_BITS'd1887992368, `RNS_PRIME_BITS'd836979688, `RNS_PRIME_BITS'd515006513, `RNS_PRIME_BITS'd1668241126, `RNS_PRIME_BITS'd2026491722, `RNS_PRIME_BITS'd2133408314, `RNS_PRIME_BITS'd989798598, `RNS_PRIME_BITS'd555817760},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd2011503780, `RNS_PRIME_BITS'd1241115807, `RNS_PRIME_BITS'd1926727251, `RNS_PRIME_BITS'd1417120048, `RNS_PRIME_BITS'd1248212236, `RNS_PRIME_BITS'd1924389879, `RNS_PRIME_BITS'd433605968, `RNS_PRIME_BITS'd1767329344, `RNS_PRIME_BITS'd1343693298, `RNS_PRIME_BITS'd1349087406}
		},
		'{
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd1905608379, `RNS_PRIME_BITS'd1170697539, `RNS_PRIME_BITS'd1389758140, `RNS_PRIME_BITS'd1606412274, `RNS_PRIME_BITS'd1057462251, `RNS_PRIME_BITS'd1743432597, `RNS_PRIME_BITS'd1265131124, `RNS_PRIME_BITS'd729269125, `RNS_PRIME_BITS'd753054750, `RNS_PRIME_BITS'd1869966969},
			'{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd709247253, `RNS_PRIME_BITS'd1959674563, `RNS_PRIME_BITS'd1149910281, `RNS_PRIME_BITS'd70923878, `RNS_PRIME_BITS'd1864899372, `RNS_PRIME_BITS'd254634607, `RNS_PRIME_BITS'd430810079, `RNS_PRIME_BITS'd1820042355, `RNS_PRIME_BITS'd228849514, `RNS_PRIME_BITS'd1560995145},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1936165201, `RNS_PRIME_BITS'd1757746099, `RNS_PRIME_BITS'd765710529, `RNS_PRIME_BITS'd731708433, `RNS_PRIME_BITS'd177823550, `RNS_PRIME_BITS'd1928984916, `RNS_PRIME_BITS'd698257183, `RNS_PRIME_BITS'd612543361, `RNS_PRIME_BITS'd100680894, `RNS_PRIME_BITS'd2069754184},
			'{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd1974918850, `RNS_PRIME_BITS'd39437613, `RNS_PRIME_BITS'd1609869490, `RNS_PRIME_BITS'd1513548799, `RNS_PRIME_BITS'd1695676616, `RNS_PRIME_BITS'd1373190017, `RNS_PRIME_BITS'd907428384, `RNS_PRIME_BITS'd1003502887, `RNS_PRIME_BITS'd399471434, `RNS_PRIME_BITS'd174773545},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd1815836891, `RNS_PRIME_BITS'd302001247, `RNS_PRIME_BITS'd883769459, `RNS_PRIME_BITS'd166271429, `RNS_PRIME_BITS'd882155119, `RNS_PRIME_BITS'd773786303, `RNS_PRIME_BITS'd1391102744, `RNS_PRIME_BITS'd1901978746, `RNS_PRIME_BITS'd458605918, `RNS_PRIME_BITS'd1841739514},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd399956847, `RNS_PRIME_BITS'd351323783, `RNS_PRIME_BITS'd1139039780, `RNS_PRIME_BITS'd1848784089, `RNS_PRIME_BITS'd1126125905, `RNS_PRIME_BITS'd1222540734, `RNS_PRIME_BITS'd2053470597, `RNS_PRIME_BITS'd629785686, `RNS_PRIME_BITS'd1241293996, `RNS_PRIME_BITS'd1520072791},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd284085739, `RNS_PRIME_BITS'd266313492, `RNS_PRIME_BITS'd2040458950, `RNS_PRIME_BITS'd310927866, `RNS_PRIME_BITS'd628013457, `RNS_PRIME_BITS'd663477868, `RNS_PRIME_BITS'd429897855, `RNS_PRIME_BITS'd1965958989, `RNS_PRIME_BITS'd1434991268, `RNS_PRIME_BITS'd1751195530},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd569519112, `RNS_PRIME_BITS'd44203046, `RNS_PRIME_BITS'd769743762, `RNS_PRIME_BITS'd1077380974, `RNS_PRIME_BITS'd1228025889, `RNS_PRIME_BITS'd1152375492, `RNS_PRIME_BITS'd1958929741, `RNS_PRIME_BITS'd312023942, `RNS_PRIME_BITS'd1474011863, `RNS_PRIME_BITS'd799660867},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd360457343, `RNS_PRIME_BITS'd20515705, `RNS_PRIME_BITS'd1280981765, `RNS_PRIME_BITS'd617710037, `RNS_PRIME_BITS'd1859265536, `RNS_PRIME_BITS'd1694423570, `RNS_PRIME_BITS'd291827467, `RNS_PRIME_BITS'd1742260953, `RNS_PRIME_BITS'd1640934552, `RNS_PRIME_BITS'd220406061},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd1166498747, `RNS_PRIME_BITS'd763502739, `RNS_PRIME_BITS'd701694283, `RNS_PRIME_BITS'd1261723735, `RNS_PRIME_BITS'd1132036341, `RNS_PRIME_BITS'd1913190995, `RNS_PRIME_BITS'd1620503003, `RNS_PRIME_BITS'd979625160, `RNS_PRIME_BITS'd2015345379, `RNS_PRIME_BITS'd324899018},
			'{`RNS_PRIME_BITS'd152, `RNS_PRIME_BITS'd1611229087, `RNS_PRIME_BITS'd455967556, `RNS_PRIME_BITS'd1412439266, `RNS_PRIME_BITS'd980326232, `RNS_PRIME_BITS'd1419341904, `RNS_PRIME_BITS'd1379750018, `RNS_PRIME_BITS'd469290645, `RNS_PRIME_BITS'd1981826023, `RNS_PRIME_BITS'd562020848, `RNS_PRIME_BITS'd1531228116},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1227167173, `RNS_PRIME_BITS'd408464823, `RNS_PRIME_BITS'd495814057, `RNS_PRIME_BITS'd889456575, `RNS_PRIME_BITS'd932180381, `RNS_PRIME_BITS'd2121582464, `RNS_PRIME_BITS'd623989577, `RNS_PRIME_BITS'd1503131402, `RNS_PRIME_BITS'd880571920, `RNS_PRIME_BITS'd708130909},
			'{`RNS_PRIME_BITS'd188, `RNS_PRIME_BITS'd1800130525, `RNS_PRIME_BITS'd834512112, `RNS_PRIME_BITS'd1503346161, `RNS_PRIME_BITS'd473295986, `RNS_PRIME_BITS'd469184641, `RNS_PRIME_BITS'd667684583, `RNS_PRIME_BITS'd358466462, `RNS_PRIME_BITS'd1792895807, `RNS_PRIME_BITS'd1413609744, `RNS_PRIME_BITS'd1935251909},
			'{`RNS_PRIME_BITS'd37, `RNS_PRIME_BITS'd1335457321, `RNS_PRIME_BITS'd2070414142, `RNS_PRIME_BITS'd1133934464, `RNS_PRIME_BITS'd1513352, `RNS_PRIME_BITS'd70870521, `RNS_PRIME_BITS'd962752820, `RNS_PRIME_BITS'd1798268636, `RNS_PRIME_BITS'd1766817016, `RNS_PRIME_BITS'd550652678, `RNS_PRIME_BITS'd1904135228},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd101758966, `RNS_PRIME_BITS'd1987927726, `RNS_PRIME_BITS'd338714856, `RNS_PRIME_BITS'd15177129, `RNS_PRIME_BITS'd2125111826, `RNS_PRIME_BITS'd1091642268, `RNS_PRIME_BITS'd2046420475, `RNS_PRIME_BITS'd35371964, `RNS_PRIME_BITS'd1709435439, `RNS_PRIME_BITS'd265583765},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1310920260, `RNS_PRIME_BITS'd687504166, `RNS_PRIME_BITS'd987937166, `RNS_PRIME_BITS'd1906589986, `RNS_PRIME_BITS'd1990591242, `RNS_PRIME_BITS'd1675370977, `RNS_PRIME_BITS'd496807822, `RNS_PRIME_BITS'd978560938, `RNS_PRIME_BITS'd173669004, `RNS_PRIME_BITS'd953490765},
			'{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd930090834, `RNS_PRIME_BITS'd2123097026, `RNS_PRIME_BITS'd412613716, `RNS_PRIME_BITS'd1031919483, `RNS_PRIME_BITS'd358153426, `RNS_PRIME_BITS'd331689246, `RNS_PRIME_BITS'd222136494, `RNS_PRIME_BITS'd1235484335, `RNS_PRIME_BITS'd1396395649, `RNS_PRIME_BITS'd469356860},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd270249878, `RNS_PRIME_BITS'd389472032, `RNS_PRIME_BITS'd1505692275, `RNS_PRIME_BITS'd440637273, `RNS_PRIME_BITS'd334302497, `RNS_PRIME_BITS'd970013484, `RNS_PRIME_BITS'd765115485, `RNS_PRIME_BITS'd1405808946, `RNS_PRIME_BITS'd1988196252, `RNS_PRIME_BITS'd814888933},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd726647235, `RNS_PRIME_BITS'd1969799553, `RNS_PRIME_BITS'd119866544, `RNS_PRIME_BITS'd1502131067, `RNS_PRIME_BITS'd387749296, `RNS_PRIME_BITS'd1567137653, `RNS_PRIME_BITS'd308762201, `RNS_PRIME_BITS'd1209995003, `RNS_PRIME_BITS'd740031860, `RNS_PRIME_BITS'd1674634276},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1611912133, `RNS_PRIME_BITS'd2095481433, `RNS_PRIME_BITS'd262813511, `RNS_PRIME_BITS'd658686310, `RNS_PRIME_BITS'd1987417067, `RNS_PRIME_BITS'd154583239, `RNS_PRIME_BITS'd1689858097, `RNS_PRIME_BITS'd359979316, `RNS_PRIME_BITS'd325314415, `RNS_PRIME_BITS'd1503495923},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd552841867, `RNS_PRIME_BITS'd393882620, `RNS_PRIME_BITS'd1667324748, `RNS_PRIME_BITS'd789366687, `RNS_PRIME_BITS'd1869073001, `RNS_PRIME_BITS'd1706227453, `RNS_PRIME_BITS'd2064059329, `RNS_PRIME_BITS'd2090703674, `RNS_PRIME_BITS'd947892668, `RNS_PRIME_BITS'd118868154},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd390596015, `RNS_PRIME_BITS'd1788869713, `RNS_PRIME_BITS'd284948187, `RNS_PRIME_BITS'd1640431632, `RNS_PRIME_BITS'd1823174010, `RNS_PRIME_BITS'd155906171, `RNS_PRIME_BITS'd2049865255, `RNS_PRIME_BITS'd455138144, `RNS_PRIME_BITS'd413929046, `RNS_PRIME_BITS'd65917259},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd912522155, `RNS_PRIME_BITS'd739704467, `RNS_PRIME_BITS'd872116099, `RNS_PRIME_BITS'd931598226, `RNS_PRIME_BITS'd1241933811, `RNS_PRIME_BITS'd1256002517, `RNS_PRIME_BITS'd323316556, `RNS_PRIME_BITS'd1684147304, `RNS_PRIME_BITS'd1584164385, `RNS_PRIME_BITS'd1334857965},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd848695442, `RNS_PRIME_BITS'd301951100, `RNS_PRIME_BITS'd1044279592, `RNS_PRIME_BITS'd825439986, `RNS_PRIME_BITS'd1598509399, `RNS_PRIME_BITS'd2129591830, `RNS_PRIME_BITS'd287659788, `RNS_PRIME_BITS'd687852664, `RNS_PRIME_BITS'd1336394461, `RNS_PRIME_BITS'd842862749},
			'{`RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd1692757107, `RNS_PRIME_BITS'd917084715, `RNS_PRIME_BITS'd420851668, `RNS_PRIME_BITS'd1954192912, `RNS_PRIME_BITS'd1465203506, `RNS_PRIME_BITS'd1924292289, `RNS_PRIME_BITS'd1912481428, `RNS_PRIME_BITS'd2016268741, `RNS_PRIME_BITS'd1235328263, `RNS_PRIME_BITS'd618866336},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd903648270, `RNS_PRIME_BITS'd174679689, `RNS_PRIME_BITS'd143897686, `RNS_PRIME_BITS'd854253824, `RNS_PRIME_BITS'd2021158380, `RNS_PRIME_BITS'd1479812437, `RNS_PRIME_BITS'd555705564, `RNS_PRIME_BITS'd1169146205, `RNS_PRIME_BITS'd296778544, `RNS_PRIME_BITS'd346506097},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd1261704741, `RNS_PRIME_BITS'd465659126, `RNS_PRIME_BITS'd280734625, `RNS_PRIME_BITS'd1294704138, `RNS_PRIME_BITS'd560141073, `RNS_PRIME_BITS'd1965990246, `RNS_PRIME_BITS'd1646233431, `RNS_PRIME_BITS'd1743286156, `RNS_PRIME_BITS'd2077586176, `RNS_PRIME_BITS'd1757906155},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd1745751452, `RNS_PRIME_BITS'd787770100, `RNS_PRIME_BITS'd1609074435, `RNS_PRIME_BITS'd908002122, `RNS_PRIME_BITS'd416136957, `RNS_PRIME_BITS'd2132813960, `RNS_PRIME_BITS'd1205370639, `RNS_PRIME_BITS'd1986777395, `RNS_PRIME_BITS'd1699089572, `RNS_PRIME_BITS'd416596136},
			'{`RNS_PRIME_BITS'd91, `RNS_PRIME_BITS'd1662489650, `RNS_PRIME_BITS'd1099040322, `RNS_PRIME_BITS'd618970414, `RNS_PRIME_BITS'd1660124537, `RNS_PRIME_BITS'd1900475151, `RNS_PRIME_BITS'd402857968, `RNS_PRIME_BITS'd1006178035, `RNS_PRIME_BITS'd957284596, `RNS_PRIME_BITS'd336255261, `RNS_PRIME_BITS'd1643280197},
			'{`RNS_PRIME_BITS'd109, `RNS_PRIME_BITS'd1190035208, `RNS_PRIME_BITS'd1516930969, `RNS_PRIME_BITS'd797448021, `RNS_PRIME_BITS'd1145485194, `RNS_PRIME_BITS'd768463650, `RNS_PRIME_BITS'd570210368, `RNS_PRIME_BITS'd1253624501, `RNS_PRIME_BITS'd994683233, `RNS_PRIME_BITS'd1775817556, `RNS_PRIME_BITS'd1210365831},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd95795481, `RNS_PRIME_BITS'd707762392, `RNS_PRIME_BITS'd1232181897, `RNS_PRIME_BITS'd1373266689, `RNS_PRIME_BITS'd948758173, `RNS_PRIME_BITS'd1381259791, `RNS_PRIME_BITS'd667074869, `RNS_PRIME_BITS'd427321030, `RNS_PRIME_BITS'd923915746, `RNS_PRIME_BITS'd22655282},
			'{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd467744686, `RNS_PRIME_BITS'd1547401623, `RNS_PRIME_BITS'd557313088, `RNS_PRIME_BITS'd20295905, `RNS_PRIME_BITS'd66217269, `RNS_PRIME_BITS'd2085233349, `RNS_PRIME_BITS'd617714744, `RNS_PRIME_BITS'd316881717, `RNS_PRIME_BITS'd75147898, `RNS_PRIME_BITS'd1629310436},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd880712458, `RNS_PRIME_BITS'd920108742, `RNS_PRIME_BITS'd2079661876, `RNS_PRIME_BITS'd1013783995, `RNS_PRIME_BITS'd895185233, `RNS_PRIME_BITS'd1189568688, `RNS_PRIME_BITS'd163112484, `RNS_PRIME_BITS'd1597079095, `RNS_PRIME_BITS'd1103395311, `RNS_PRIME_BITS'd1698428070},
			'{`RNS_PRIME_BITS'd170, `RNS_PRIME_BITS'd1033605430, `RNS_PRIME_BITS'd886085760, `RNS_PRIME_BITS'd1223225088, `RNS_PRIME_BITS'd897292109, `RNS_PRIME_BITS'd311997283, `RNS_PRIME_BITS'd258735397, `RNS_PRIME_BITS'd812053791, `RNS_PRIME_BITS'd986488792, `RNS_PRIME_BITS'd1881406373, `RNS_PRIME_BITS'd1078738177},
			'{`RNS_PRIME_BITS'd196, `RNS_PRIME_BITS'd320038852, `RNS_PRIME_BITS'd1863324439, `RNS_PRIME_BITS'd452315465, `RNS_PRIME_BITS'd1334095, `RNS_PRIME_BITS'd2047712474, `RNS_PRIME_BITS'd855657194, `RNS_PRIME_BITS'd906932808, `RNS_PRIME_BITS'd1010280612, `RNS_PRIME_BITS'd52786527, `RNS_PRIME_BITS'd1548651225},
			'{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd1796187890, `RNS_PRIME_BITS'd1952376485, `RNS_PRIME_BITS'd767184907, `RNS_PRIME_BITS'd597049005, `RNS_PRIME_BITS'd1757755239, `RNS_PRIME_BITS'd105918204, `RNS_PRIME_BITS'd508880001, `RNS_PRIME_BITS'd842657938, `RNS_PRIME_BITS'd2028506104, `RNS_PRIME_BITS'd1919617695},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd377765506, `RNS_PRIME_BITS'd1533466317, `RNS_PRIME_BITS'd997783072, `RNS_PRIME_BITS'd66563855, `RNS_PRIME_BITS'd484254400, `RNS_PRIME_BITS'd298474816, `RNS_PRIME_BITS'd445692858, `RNS_PRIME_BITS'd321770165, `RNS_PRIME_BITS'd1208725747, `RNS_PRIME_BITS'd925170256},
			'{`RNS_PRIME_BITS'd180, `RNS_PRIME_BITS'd2126785476, `RNS_PRIME_BITS'd1367193419, `RNS_PRIME_BITS'd545731695, `RNS_PRIME_BITS'd1387825439, `RNS_PRIME_BITS'd582312990, `RNS_PRIME_BITS'd1582369776, `RNS_PRIME_BITS'd666646831, `RNS_PRIME_BITS'd1365996028, `RNS_PRIME_BITS'd2095999815, `RNS_PRIME_BITS'd719915030},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd834118430, `RNS_PRIME_BITS'd1435998463, `RNS_PRIME_BITS'd2092360347, `RNS_PRIME_BITS'd2117517657, `RNS_PRIME_BITS'd260510533, `RNS_PRIME_BITS'd1930785237, `RNS_PRIME_BITS'd1703467625, `RNS_PRIME_BITS'd165336970, `RNS_PRIME_BITS'd839521087, `RNS_PRIME_BITS'd1526137028},
			'{`RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd1051425869, `RNS_PRIME_BITS'd415623283, `RNS_PRIME_BITS'd2048635488, `RNS_PRIME_BITS'd1056331181, `RNS_PRIME_BITS'd514754326, `RNS_PRIME_BITS'd218175788, `RNS_PRIME_BITS'd1489271734, `RNS_PRIME_BITS'd167900506, `RNS_PRIME_BITS'd2103010075, `RNS_PRIME_BITS'd179162060},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd1963006511, `RNS_PRIME_BITS'd468087279, `RNS_PRIME_BITS'd1651996066, `RNS_PRIME_BITS'd1088493537, `RNS_PRIME_BITS'd1405533987, `RNS_PRIME_BITS'd1700050967, `RNS_PRIME_BITS'd2063895364, `RNS_PRIME_BITS'd318579839, `RNS_PRIME_BITS'd30697162, `RNS_PRIME_BITS'd65880226},
			'{`RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd702756135, `RNS_PRIME_BITS'd1007328570, `RNS_PRIME_BITS'd1922822338, `RNS_PRIME_BITS'd1966632641, `RNS_PRIME_BITS'd1858307026, `RNS_PRIME_BITS'd1436162338, `RNS_PRIME_BITS'd275116871, `RNS_PRIME_BITS'd1612436804, `RNS_PRIME_BITS'd1891753254, `RNS_PRIME_BITS'd1868195849},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd817496138, `RNS_PRIME_BITS'd338330661, `RNS_PRIME_BITS'd1888054724, `RNS_PRIME_BITS'd1421952796, `RNS_PRIME_BITS'd2123423669, `RNS_PRIME_BITS'd1790144218, `RNS_PRIME_BITS'd1628337834, `RNS_PRIME_BITS'd1961413114, `RNS_PRIME_BITS'd992822690, `RNS_PRIME_BITS'd942331185},
			'{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd1171275869, `RNS_PRIME_BITS'd720470275, `RNS_PRIME_BITS'd1715851322, `RNS_PRIME_BITS'd65145786, `RNS_PRIME_BITS'd1692006233, `RNS_PRIME_BITS'd1961168146, `RNS_PRIME_BITS'd453261293, `RNS_PRIME_BITS'd690505322, `RNS_PRIME_BITS'd1729084170, `RNS_PRIME_BITS'd685584863},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd237031139, `RNS_PRIME_BITS'd332724881, `RNS_PRIME_BITS'd297337988, `RNS_PRIME_BITS'd1741706420, `RNS_PRIME_BITS'd1103181801, `RNS_PRIME_BITS'd54349747, `RNS_PRIME_BITS'd1601488263, `RNS_PRIME_BITS'd1473433585, `RNS_PRIME_BITS'd1668060765, `RNS_PRIME_BITS'd826559556},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd1128970952, `RNS_PRIME_BITS'd743687105, `RNS_PRIME_BITS'd915545864, `RNS_PRIME_BITS'd1049117552, `RNS_PRIME_BITS'd1263680574, `RNS_PRIME_BITS'd251419754, `RNS_PRIME_BITS'd1809744746, `RNS_PRIME_BITS'd1930328758, `RNS_PRIME_BITS'd1558662361, `RNS_PRIME_BITS'd1423892144},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd2066884645, `RNS_PRIME_BITS'd1802028247, `RNS_PRIME_BITS'd52102155, `RNS_PRIME_BITS'd480998964, `RNS_PRIME_BITS'd738884885, `RNS_PRIME_BITS'd357172811, `RNS_PRIME_BITS'd1096125755, `RNS_PRIME_BITS'd418510638, `RNS_PRIME_BITS'd448191408, `RNS_PRIME_BITS'd624764735},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd364130156, `RNS_PRIME_BITS'd1814992890, `RNS_PRIME_BITS'd1456610446, `RNS_PRIME_BITS'd519575641, `RNS_PRIME_BITS'd1454843701, `RNS_PRIME_BITS'd1029398513, `RNS_PRIME_BITS'd1033443501, `RNS_PRIME_BITS'd942739069, `RNS_PRIME_BITS'd946512577, `RNS_PRIME_BITS'd1315660026},
			'{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd1845704137, `RNS_PRIME_BITS'd1460160736, `RNS_PRIME_BITS'd1578808907, `RNS_PRIME_BITS'd254551637, `RNS_PRIME_BITS'd2048044387, `RNS_PRIME_BITS'd2032254360, `RNS_PRIME_BITS'd1163608180, `RNS_PRIME_BITS'd1394982888, `RNS_PRIME_BITS'd1223825108, `RNS_PRIME_BITS'd2038500193},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd435888803, `RNS_PRIME_BITS'd988002405, `RNS_PRIME_BITS'd845883156, `RNS_PRIME_BITS'd1954048083, `RNS_PRIME_BITS'd1913232785, `RNS_PRIME_BITS'd1302560458, `RNS_PRIME_BITS'd2075998619, `RNS_PRIME_BITS'd1157659084, `RNS_PRIME_BITS'd1965853377, `RNS_PRIME_BITS'd1421494764},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1005613900, `RNS_PRIME_BITS'd1978333843, `RNS_PRIME_BITS'd504043456, `RNS_PRIME_BITS'd594762138, `RNS_PRIME_BITS'd1565374703, `RNS_PRIME_BITS'd1803362272, `RNS_PRIME_BITS'd1247581086, `RNS_PRIME_BITS'd1727361149, `RNS_PRIME_BITS'd536271744, `RNS_PRIME_BITS'd125520790},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd1481222563, `RNS_PRIME_BITS'd1855234899, `RNS_PRIME_BITS'd199836192, `RNS_PRIME_BITS'd308970543, `RNS_PRIME_BITS'd530414172, `RNS_PRIME_BITS'd627913734, `RNS_PRIME_BITS'd2143596166, `RNS_PRIME_BITS'd1206180128, `RNS_PRIME_BITS'd1332288065, `RNS_PRIME_BITS'd972389562},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd559220682, `RNS_PRIME_BITS'd1046244715, `RNS_PRIME_BITS'd93788787, `RNS_PRIME_BITS'd2029592528, `RNS_PRIME_BITS'd297260250, `RNS_PRIME_BITS'd431155812, `RNS_PRIME_BITS'd1465701889, `RNS_PRIME_BITS'd366486222, `RNS_PRIME_BITS'd322554010, `RNS_PRIME_BITS'd1922559236},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd879038792, `RNS_PRIME_BITS'd2121109936, `RNS_PRIME_BITS'd2101922480, `RNS_PRIME_BITS'd1501566639, `RNS_PRIME_BITS'd2060965004, `RNS_PRIME_BITS'd662200455, `RNS_PRIME_BITS'd1865759069, `RNS_PRIME_BITS'd1733380592, `RNS_PRIME_BITS'd210083102, `RNS_PRIME_BITS'd1004150580},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd1500423343, `RNS_PRIME_BITS'd94385508, `RNS_PRIME_BITS'd344041825, `RNS_PRIME_BITS'd723054482, `RNS_PRIME_BITS'd1297453453, `RNS_PRIME_BITS'd41488238, `RNS_PRIME_BITS'd1462067684, `RNS_PRIME_BITS'd1960502620, `RNS_PRIME_BITS'd2086988844, `RNS_PRIME_BITS'd1214499461},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd2083574133, `RNS_PRIME_BITS'd829976384, `RNS_PRIME_BITS'd189978152, `RNS_PRIME_BITS'd2045744174, `RNS_PRIME_BITS'd1720705220, `RNS_PRIME_BITS'd505021027, `RNS_PRIME_BITS'd184462552, `RNS_PRIME_BITS'd1401715667, `RNS_PRIME_BITS'd829160128, `RNS_PRIME_BITS'd904612413},
			'{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd1209403816, `RNS_PRIME_BITS'd586389397, `RNS_PRIME_BITS'd1921920701, `RNS_PRIME_BITS'd299152541, `RNS_PRIME_BITS'd745941080, `RNS_PRIME_BITS'd439025579, `RNS_PRIME_BITS'd638729448, `RNS_PRIME_BITS'd2119618454, `RNS_PRIME_BITS'd1697564957, `RNS_PRIME_BITS'd1760568699},
			'{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd678620432, `RNS_PRIME_BITS'd933085404, `RNS_PRIME_BITS'd815336414, `RNS_PRIME_BITS'd1742297440, `RNS_PRIME_BITS'd1733176698, `RNS_PRIME_BITS'd250893959, `RNS_PRIME_BITS'd1728841612, `RNS_PRIME_BITS'd196185798, `RNS_PRIME_BITS'd1522287068, `RNS_PRIME_BITS'd1302305588},
			'{`RNS_PRIME_BITS'd140, `RNS_PRIME_BITS'd881599791, `RNS_PRIME_BITS'd217582950, `RNS_PRIME_BITS'd1199221674, `RNS_PRIME_BITS'd1228275556, `RNS_PRIME_BITS'd2056883187, `RNS_PRIME_BITS'd1336084535, `RNS_PRIME_BITS'd1372314211, `RNS_PRIME_BITS'd124585053, `RNS_PRIME_BITS'd865467042, `RNS_PRIME_BITS'd1913363758},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd2044793122, `RNS_PRIME_BITS'd411601935, `RNS_PRIME_BITS'd124780452, `RNS_PRIME_BITS'd731200665, `RNS_PRIME_BITS'd1017329313, `RNS_PRIME_BITS'd692806430, `RNS_PRIME_BITS'd531360161, `RNS_PRIME_BITS'd1804011624, `RNS_PRIME_BITS'd949932524, `RNS_PRIME_BITS'd1764124780},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd2084397288, `RNS_PRIME_BITS'd961515945, `RNS_PRIME_BITS'd2007610731, `RNS_PRIME_BITS'd2115985192, `RNS_PRIME_BITS'd931598540, `RNS_PRIME_BITS'd698432291, `RNS_PRIME_BITS'd2122069994, `RNS_PRIME_BITS'd2059347814, `RNS_PRIME_BITS'd918764298, `RNS_PRIME_BITS'd1126086117},
			'{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd400869838, `RNS_PRIME_BITS'd75154276, `RNS_PRIME_BITS'd1852773008, `RNS_PRIME_BITS'd1458042808, `RNS_PRIME_BITS'd669713673, `RNS_PRIME_BITS'd1510460000, `RNS_PRIME_BITS'd1822636613, `RNS_PRIME_BITS'd1512813193, `RNS_PRIME_BITS'd1194372006, `RNS_PRIME_BITS'd1093745618},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd1348413174, `RNS_PRIME_BITS'd1343161778, `RNS_PRIME_BITS'd399981772, `RNS_PRIME_BITS'd1168193404, `RNS_PRIME_BITS'd1835663555, `RNS_PRIME_BITS'd556489014, `RNS_PRIME_BITS'd1143521926, `RNS_PRIME_BITS'd1450703842, `RNS_PRIME_BITS'd814204318, `RNS_PRIME_BITS'd1085380418},
			'{`RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd1455949476, `RNS_PRIME_BITS'd997202604, `RNS_PRIME_BITS'd1253597608, `RNS_PRIME_BITS'd1867996744, `RNS_PRIME_BITS'd475684206, `RNS_PRIME_BITS'd689847630, `RNS_PRIME_BITS'd1645440166, `RNS_PRIME_BITS'd899610637, `RNS_PRIME_BITS'd99936376, `RNS_PRIME_BITS'd1769166010}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd2057247496, `RNS_PRIME_BITS'd779215751, `RNS_PRIME_BITS'd370435910, `RNS_PRIME_BITS'd841973641, `RNS_PRIME_BITS'd475364771, `RNS_PRIME_BITS'd231690204, `RNS_PRIME_BITS'd1541415722, `RNS_PRIME_BITS'd194871934, `RNS_PRIME_BITS'd886072123, `RNS_PRIME_BITS'd1865704193},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd1260554722, `RNS_PRIME_BITS'd1686205273, `RNS_PRIME_BITS'd1676246087, `RNS_PRIME_BITS'd601725004, `RNS_PRIME_BITS'd1052990186, `RNS_PRIME_BITS'd1780898339, `RNS_PRIME_BITS'd1659717421, `RNS_PRIME_BITS'd1213377041, `RNS_PRIME_BITS'd1443647279, `RNS_PRIME_BITS'd1754929589},
			'{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd10246935, `RNS_PRIME_BITS'd636930725, `RNS_PRIME_BITS'd1155520764, `RNS_PRIME_BITS'd618280203, `RNS_PRIME_BITS'd1782162664, `RNS_PRIME_BITS'd695430977, `RNS_PRIME_BITS'd454849180, `RNS_PRIME_BITS'd614591563, `RNS_PRIME_BITS'd1702422973, `RNS_PRIME_BITS'd1980125346},
			'{`RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd266682724, `RNS_PRIME_BITS'd854529560, `RNS_PRIME_BITS'd1652445821, `RNS_PRIME_BITS'd1234313022, `RNS_PRIME_BITS'd730731559, `RNS_PRIME_BITS'd1171413732, `RNS_PRIME_BITS'd295262243, `RNS_PRIME_BITS'd625585397, `RNS_PRIME_BITS'd1312322519, `RNS_PRIME_BITS'd796672691},
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd944093942, `RNS_PRIME_BITS'd18818776, `RNS_PRIME_BITS'd1171301610, `RNS_PRIME_BITS'd453102958, `RNS_PRIME_BITS'd718126580, `RNS_PRIME_BITS'd2133126524, `RNS_PRIME_BITS'd1635475949, `RNS_PRIME_BITS'd435243418, `RNS_PRIME_BITS'd403897523, `RNS_PRIME_BITS'd1200997362},
			'{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd231350874, `RNS_PRIME_BITS'd472445870, `RNS_PRIME_BITS'd1987717261, `RNS_PRIME_BITS'd1256235188, `RNS_PRIME_BITS'd2145048151, `RNS_PRIME_BITS'd685077107, `RNS_PRIME_BITS'd1463158621, `RNS_PRIME_BITS'd10698702, `RNS_PRIME_BITS'd457606687, `RNS_PRIME_BITS'd902646604},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd204955343, `RNS_PRIME_BITS'd1375940579, `RNS_PRIME_BITS'd1695452320, `RNS_PRIME_BITS'd253932424, `RNS_PRIME_BITS'd1688282148, `RNS_PRIME_BITS'd120353182, `RNS_PRIME_BITS'd1445378361, `RNS_PRIME_BITS'd1942196180, `RNS_PRIME_BITS'd709506112, `RNS_PRIME_BITS'd784521215},
			'{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd1851001298, `RNS_PRIME_BITS'd1368164498, `RNS_PRIME_BITS'd1410975001, `RNS_PRIME_BITS'd30385488, `RNS_PRIME_BITS'd922712315, `RNS_PRIME_BITS'd550224444, `RNS_PRIME_BITS'd1284005195, `RNS_PRIME_BITS'd1992318958, `RNS_PRIME_BITS'd1565077607, `RNS_PRIME_BITS'd742563801},
			'{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd1841082732, `RNS_PRIME_BITS'd324630693, `RNS_PRIME_BITS'd1228850860, `RNS_PRIME_BITS'd1326469721, `RNS_PRIME_BITS'd141710441, `RNS_PRIME_BITS'd380169378, `RNS_PRIME_BITS'd1003363831, `RNS_PRIME_BITS'd396925408, `RNS_PRIME_BITS'd856738281, `RNS_PRIME_BITS'd13355984},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1695631662, `RNS_PRIME_BITS'd1112453373, `RNS_PRIME_BITS'd78575208, `RNS_PRIME_BITS'd2130972150, `RNS_PRIME_BITS'd2108004692, `RNS_PRIME_BITS'd1363733948, `RNS_PRIME_BITS'd858064176, `RNS_PRIME_BITS'd1393568189, `RNS_PRIME_BITS'd388160252, `RNS_PRIME_BITS'd599942071},
			'{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd417142305, `RNS_PRIME_BITS'd800749392, `RNS_PRIME_BITS'd198746382, `RNS_PRIME_BITS'd4114996, `RNS_PRIME_BITS'd1198663949, `RNS_PRIME_BITS'd1097586735, `RNS_PRIME_BITS'd831202174, `RNS_PRIME_BITS'd351639504, `RNS_PRIME_BITS'd742809771, `RNS_PRIME_BITS'd1974434026},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd1663061988, `RNS_PRIME_BITS'd1383427189, `RNS_PRIME_BITS'd946179966, `RNS_PRIME_BITS'd1014462323, `RNS_PRIME_BITS'd223127606, `RNS_PRIME_BITS'd633006660, `RNS_PRIME_BITS'd1601845436, `RNS_PRIME_BITS'd1754522162, `RNS_PRIME_BITS'd1898410778, `RNS_PRIME_BITS'd654113139},
			'{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd965437543, `RNS_PRIME_BITS'd887691573, `RNS_PRIME_BITS'd1792110841, `RNS_PRIME_BITS'd1617361755, `RNS_PRIME_BITS'd834751540, `RNS_PRIME_BITS'd1778860263, `RNS_PRIME_BITS'd1569099260, `RNS_PRIME_BITS'd823497743, `RNS_PRIME_BITS'd1743674651, `RNS_PRIME_BITS'd1901036331},
			'{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd1864304537, `RNS_PRIME_BITS'd324956842, `RNS_PRIME_BITS'd1860432042, `RNS_PRIME_BITS'd610330943, `RNS_PRIME_BITS'd1827026737, `RNS_PRIME_BITS'd876332408, `RNS_PRIME_BITS'd832568892, `RNS_PRIME_BITS'd2046806424, `RNS_PRIME_BITS'd1553373517, `RNS_PRIME_BITS'd780926028},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd468548188, `RNS_PRIME_BITS'd1314765770, `RNS_PRIME_BITS'd504576663, `RNS_PRIME_BITS'd113932602, `RNS_PRIME_BITS'd860852631, `RNS_PRIME_BITS'd171226679, `RNS_PRIME_BITS'd1157748724, `RNS_PRIME_BITS'd530530516, `RNS_PRIME_BITS'd373438624, `RNS_PRIME_BITS'd394397221},
			'{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd773682191, `RNS_PRIME_BITS'd1969063420, `RNS_PRIME_BITS'd596897602, `RNS_PRIME_BITS'd1584589556, `RNS_PRIME_BITS'd543805312, `RNS_PRIME_BITS'd833826561, `RNS_PRIME_BITS'd1136182139, `RNS_PRIME_BITS'd167251796, `RNS_PRIME_BITS'd705767662, `RNS_PRIME_BITS'd2110628826},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd730823491, `RNS_PRIME_BITS'd1498044159, `RNS_PRIME_BITS'd1103805929, `RNS_PRIME_BITS'd1796874967, `RNS_PRIME_BITS'd2055014391, `RNS_PRIME_BITS'd738216900, `RNS_PRIME_BITS'd22555559, `RNS_PRIME_BITS'd1331147409, `RNS_PRIME_BITS'd169450983, `RNS_PRIME_BITS'd857406704},
			'{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd2040069578, `RNS_PRIME_BITS'd1588951895, `RNS_PRIME_BITS'd1231303236, `RNS_PRIME_BITS'd106480088, `RNS_PRIME_BITS'd1430130807, `RNS_PRIME_BITS'd1359112323, `RNS_PRIME_BITS'd1519108459, `RNS_PRIME_BITS'd1790981620, `RNS_PRIME_BITS'd1676746852, `RNS_PRIME_BITS'd2084063874},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd1525495041, `RNS_PRIME_BITS'd545306760, `RNS_PRIME_BITS'd2049642140, `RNS_PRIME_BITS'd1518081159, `RNS_PRIME_BITS'd1870516872, `RNS_PRIME_BITS'd644316462, `RNS_PRIME_BITS'd1837187963, `RNS_PRIME_BITS'd745292117, `RNS_PRIME_BITS'd489980081, `RNS_PRIME_BITS'd202252850},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd1467649310, `RNS_PRIME_BITS'd712277609, `RNS_PRIME_BITS'd227600337, `RNS_PRIME_BITS'd1166954678, `RNS_PRIME_BITS'd1708585294, `RNS_PRIME_BITS'd871651933, `RNS_PRIME_BITS'd864417503, `RNS_PRIME_BITS'd174379735, `RNS_PRIME_BITS'd545402836, `RNS_PRIME_BITS'd1493867213},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd642055425, `RNS_PRIME_BITS'd1634504124, `RNS_PRIME_BITS'd475255818, `RNS_PRIME_BITS'd756043802, `RNS_PRIME_BITS'd180825194, `RNS_PRIME_BITS'd623313599, `RNS_PRIME_BITS'd227633492, `RNS_PRIME_BITS'd685983244, `RNS_PRIME_BITS'd185410488, `RNS_PRIME_BITS'd753935864},
			'{`RNS_PRIME_BITS'd170, `RNS_PRIME_BITS'd1484824032, `RNS_PRIME_BITS'd1922392897, `RNS_PRIME_BITS'd893423601, `RNS_PRIME_BITS'd1745766589, `RNS_PRIME_BITS'd1196927437, `RNS_PRIME_BITS'd1212069880, `RNS_PRIME_BITS'd1920096125, `RNS_PRIME_BITS'd785824837, `RNS_PRIME_BITS'd1395293070, `RNS_PRIME_BITS'd183262496},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1310571091, `RNS_PRIME_BITS'd98277484, `RNS_PRIME_BITS'd1149083269, `RNS_PRIME_BITS'd1289949497, `RNS_PRIME_BITS'd407114305, `RNS_PRIME_BITS'd2015563283, `RNS_PRIME_BITS'd1948436391, `RNS_PRIME_BITS'd125077476, `RNS_PRIME_BITS'd1180053466, `RNS_PRIME_BITS'd2089060444},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1764811523, `RNS_PRIME_BITS'd799073470, `RNS_PRIME_BITS'd775947845, `RNS_PRIME_BITS'd2044095967, `RNS_PRIME_BITS'd2099739143, `RNS_PRIME_BITS'd295990995, `RNS_PRIME_BITS'd584899662, `RNS_PRIME_BITS'd996536362, `RNS_PRIME_BITS'd1306341838, `RNS_PRIME_BITS'd1102548026},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd124594465, `RNS_PRIME_BITS'd1618203156, `RNS_PRIME_BITS'd2029612303, `RNS_PRIME_BITS'd684986915, `RNS_PRIME_BITS'd342251377, `RNS_PRIME_BITS'd1616937730, `RNS_PRIME_BITS'd1153924893, `RNS_PRIME_BITS'd90626268, `RNS_PRIME_BITS'd691759787, `RNS_PRIME_BITS'd567705536},
			'{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd1451709026, `RNS_PRIME_BITS'd1188248873, `RNS_PRIME_BITS'd1358291083, `RNS_PRIME_BITS'd859443043, `RNS_PRIME_BITS'd1816038672, `RNS_PRIME_BITS'd1336442345, `RNS_PRIME_BITS'd988534829, `RNS_PRIME_BITS'd2113210169, `RNS_PRIME_BITS'd670154973, `RNS_PRIME_BITS'd194984665},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd1886262173, `RNS_PRIME_BITS'd1671029714, `RNS_PRIME_BITS'd499231679, `RNS_PRIME_BITS'd1010222329, `RNS_PRIME_BITS'd1141231053, `RNS_PRIME_BITS'd575758966, `RNS_PRIME_BITS'd1804276355, `RNS_PRIME_BITS'd512159432, `RNS_PRIME_BITS'd1757409767, `RNS_PRIME_BITS'd952029489},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1880915214, `RNS_PRIME_BITS'd1197202320, `RNS_PRIME_BITS'd1590053241, `RNS_PRIME_BITS'd1094141467, `RNS_PRIME_BITS'd2125381429, `RNS_PRIME_BITS'd1770765532, `RNS_PRIME_BITS'd1203644095, `RNS_PRIME_BITS'd93460477, `RNS_PRIME_BITS'd869392673, `RNS_PRIME_BITS'd1481708585},
			'{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd258040899, `RNS_PRIME_BITS'd785144572, `RNS_PRIME_BITS'd645761479, `RNS_PRIME_BITS'd1517514677, `RNS_PRIME_BITS'd1308306878, `RNS_PRIME_BITS'd1390879030, `RNS_PRIME_BITS'd1981744159, `RNS_PRIME_BITS'd696043315, `RNS_PRIME_BITS'd1382665519, `RNS_PRIME_BITS'd62593562},
			'{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd1233238386, `RNS_PRIME_BITS'd489772901, `RNS_PRIME_BITS'd1311040903, `RNS_PRIME_BITS'd1513710410, `RNS_PRIME_BITS'd285688971, `RNS_PRIME_BITS'd1697715535, `RNS_PRIME_BITS'd1390118221, `RNS_PRIME_BITS'd775519908, `RNS_PRIME_BITS'd1387084962, `RNS_PRIME_BITS'd654672642},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd571666102, `RNS_PRIME_BITS'd2092483493, `RNS_PRIME_BITS'd1553190634, `RNS_PRIME_BITS'd1052688354, `RNS_PRIME_BITS'd414052875, `RNS_PRIME_BITS'd629367403, `RNS_PRIME_BITS'd821796326, `RNS_PRIME_BITS'd1636096842, `RNS_PRIME_BITS'd1015784833, `RNS_PRIME_BITS'd447630042},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd384915487, `RNS_PRIME_BITS'd853388679, `RNS_PRIME_BITS'd840975277, `RNS_PRIME_BITS'd17174077, `RNS_PRIME_BITS'd833625985, `RNS_PRIME_BITS'd1921733263, `RNS_PRIME_BITS'd980568894, `RNS_PRIME_BITS'd25873637, `RNS_PRIME_BITS'd1359563401, `RNS_PRIME_BITS'd1927569471},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd865464910, `RNS_PRIME_BITS'd1367672206, `RNS_PRIME_BITS'd609614579, `RNS_PRIME_BITS'd486532349, `RNS_PRIME_BITS'd1628913899, `RNS_PRIME_BITS'd1991402064, `RNS_PRIME_BITS'd777005264, `RNS_PRIME_BITS'd150919199, `RNS_PRIME_BITS'd1559578338, `RNS_PRIME_BITS'd263937183},
			'{`RNS_PRIME_BITS'd91, `RNS_PRIME_BITS'd585703076, `RNS_PRIME_BITS'd245760992, `RNS_PRIME_BITS'd4306352, `RNS_PRIME_BITS'd1948360383, `RNS_PRIME_BITS'd227834606, `RNS_PRIME_BITS'd1933002616, `RNS_PRIME_BITS'd1346485866, `RNS_PRIME_BITS'd1831752628, `RNS_PRIME_BITS'd1151057459, `RNS_PRIME_BITS'd1797876074},
			'{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd460431075, `RNS_PRIME_BITS'd203171852, `RNS_PRIME_BITS'd906280681, `RNS_PRIME_BITS'd1867372021, `RNS_PRIME_BITS'd2015064892, `RNS_PRIME_BITS'd1024960624, `RNS_PRIME_BITS'd2056550803, `RNS_PRIME_BITS'd462997793, `RNS_PRIME_BITS'd1214745376, `RNS_PRIME_BITS'd1181490214},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1228367941, `RNS_PRIME_BITS'd1623532264, `RNS_PRIME_BITS'd1011352944, `RNS_PRIME_BITS'd1255071962, `RNS_PRIME_BITS'd2008770869, `RNS_PRIME_BITS'd1561013760, `RNS_PRIME_BITS'd1985013478, `RNS_PRIME_BITS'd1230926820, `RNS_PRIME_BITS'd1652167871, `RNS_PRIME_BITS'd1636931776},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd659234365, `RNS_PRIME_BITS'd2075959244, `RNS_PRIME_BITS'd1922449396, `RNS_PRIME_BITS'd1869706354, `RNS_PRIME_BITS'd1318771859, `RNS_PRIME_BITS'd1642461727, `RNS_PRIME_BITS'd891547552, `RNS_PRIME_BITS'd1395842835, `RNS_PRIME_BITS'd1332325270, `RNS_PRIME_BITS'd326002690},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd343254963, `RNS_PRIME_BITS'd2002118265, `RNS_PRIME_BITS'd879540194, `RNS_PRIME_BITS'd1042505667, `RNS_PRIME_BITS'd1864132475, `RNS_PRIME_BITS'd1070199391, `RNS_PRIME_BITS'd216215789, `RNS_PRIME_BITS'd662671173, `RNS_PRIME_BITS'd912960142, `RNS_PRIME_BITS'd1802144360},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd1591936138, `RNS_PRIME_BITS'd167015659, `RNS_PRIME_BITS'd14946662, `RNS_PRIME_BITS'd1598124643, `RNS_PRIME_BITS'd1135261976, `RNS_PRIME_BITS'd1957851369, `RNS_PRIME_BITS'd237945384, `RNS_PRIME_BITS'd244141782, `RNS_PRIME_BITS'd1746649556, `RNS_PRIME_BITS'd95627782},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd1767517112, `RNS_PRIME_BITS'd696314270, `RNS_PRIME_BITS'd1688488680, `RNS_PRIME_BITS'd1670788602, `RNS_PRIME_BITS'd154727511, `RNS_PRIME_BITS'd1614842423, `RNS_PRIME_BITS'd237735707, `RNS_PRIME_BITS'd866797377, `RNS_PRIME_BITS'd137065099, `RNS_PRIME_BITS'd784671382},
			'{`RNS_PRIME_BITS'd156, `RNS_PRIME_BITS'd717284442, `RNS_PRIME_BITS'd81389933, `RNS_PRIME_BITS'd1884303333, `RNS_PRIME_BITS'd798072551, `RNS_PRIME_BITS'd410685333, `RNS_PRIME_BITS'd1978723153, `RNS_PRIME_BITS'd1431673459, `RNS_PRIME_BITS'd12977509, `RNS_PRIME_BITS'd1034760578, `RNS_PRIME_BITS'd1140666866},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1128060383, `RNS_PRIME_BITS'd258745809, `RNS_PRIME_BITS'd1911179398, `RNS_PRIME_BITS'd1702664523, `RNS_PRIME_BITS'd2130932981, `RNS_PRIME_BITS'd382046043, `RNS_PRIME_BITS'd1129212968, `RNS_PRIME_BITS'd742974501, `RNS_PRIME_BITS'd1162158604, `RNS_PRIME_BITS'd1962492666},
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1364321915, `RNS_PRIME_BITS'd623230438, `RNS_PRIME_BITS'd353117268, `RNS_PRIME_BITS'd1783049221, `RNS_PRIME_BITS'd3315797, `RNS_PRIME_BITS'd763644073, `RNS_PRIME_BITS'd1593797503, `RNS_PRIME_BITS'd1330590062, `RNS_PRIME_BITS'd242467092, `RNS_PRIME_BITS'd240417554},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd766012726, `RNS_PRIME_BITS'd1373738953, `RNS_PRIME_BITS'd650801459, `RNS_PRIME_BITS'd372554098, `RNS_PRIME_BITS'd1540287428, `RNS_PRIME_BITS'd522940669, `RNS_PRIME_BITS'd615895277, `RNS_PRIME_BITS'd1102312905, `RNS_PRIME_BITS'd7887565, `RNS_PRIME_BITS'd1964222422},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd305896601, `RNS_PRIME_BITS'd1047035002, `RNS_PRIME_BITS'd1393401787, `RNS_PRIME_BITS'd1904778460, `RNS_PRIME_BITS'd1511043463, `RNS_PRIME_BITS'd337286337, `RNS_PRIME_BITS'd69613055, `RNS_PRIME_BITS'd1056232499, `RNS_PRIME_BITS'd521239936, `RNS_PRIME_BITS'd1989289446},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd293702305, `RNS_PRIME_BITS'd213417202, `RNS_PRIME_BITS'd1650564287, `RNS_PRIME_BITS'd1341096081, `RNS_PRIME_BITS'd1357187354, `RNS_PRIME_BITS'd778371788, `RNS_PRIME_BITS'd30696430, `RNS_PRIME_BITS'd71568482, `RNS_PRIME_BITS'd1084894881, `RNS_PRIME_BITS'd1963860413},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd2011558589, `RNS_PRIME_BITS'd209888240, `RNS_PRIME_BITS'd1730060412, `RNS_PRIME_BITS'd1531982288, `RNS_PRIME_BITS'd66160713, `RNS_PRIME_BITS'd198020266, `RNS_PRIME_BITS'd567247387, `RNS_PRIME_BITS'd1432790942, `RNS_PRIME_BITS'd2010197003, `RNS_PRIME_BITS'd699859459},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd197474236, `RNS_PRIME_BITS'd280307795, `RNS_PRIME_BITS'd131762713, `RNS_PRIME_BITS'd505826328, `RNS_PRIME_BITS'd398005689, `RNS_PRIME_BITS'd1914323495, `RNS_PRIME_BITS'd2137507732, `RNS_PRIME_BITS'd795074382, `RNS_PRIME_BITS'd1633984136, `RNS_PRIME_BITS'd144058157},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd2095984830, `RNS_PRIME_BITS'd206740997, `RNS_PRIME_BITS'd685704724, `RNS_PRIME_BITS'd505602862, `RNS_PRIME_BITS'd642488593, `RNS_PRIME_BITS'd1052124093, `RNS_PRIME_BITS'd1278494675, `RNS_PRIME_BITS'd592016439, `RNS_PRIME_BITS'd499454102, `RNS_PRIME_BITS'd281822712},
			'{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd864410747, `RNS_PRIME_BITS'd954987029, `RNS_PRIME_BITS'd1313653179, `RNS_PRIME_BITS'd1734769529, `RNS_PRIME_BITS'd2066668496, `RNS_PRIME_BITS'd937099005, `RNS_PRIME_BITS'd887790328, `RNS_PRIME_BITS'd1464077201, `RNS_PRIME_BITS'd204013155, `RNS_PRIME_BITS'd63642504},
			'{`RNS_PRIME_BITS'd101, `RNS_PRIME_BITS'd1342395238, `RNS_PRIME_BITS'd456843924, `RNS_PRIME_BITS'd1965890547, `RNS_PRIME_BITS'd1674594760, `RNS_PRIME_BITS'd224598826, `RNS_PRIME_BITS'd390738880, `RNS_PRIME_BITS'd1877793903, `RNS_PRIME_BITS'd609245160, `RNS_PRIME_BITS'd823073453, `RNS_PRIME_BITS'd1776871002},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1744489265, `RNS_PRIME_BITS'd320476356, `RNS_PRIME_BITS'd1358488152, `RNS_PRIME_BITS'd1691895170, `RNS_PRIME_BITS'd1690183888, `RNS_PRIME_BITS'd1936825693, `RNS_PRIME_BITS'd2087788190, `RNS_PRIME_BITS'd110884203, `RNS_PRIME_BITS'd333749869, `RNS_PRIME_BITS'd1637682738},
			'{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd1727982933, `RNS_PRIME_BITS'd1891498467, `RNS_PRIME_BITS'd953431164, `RNS_PRIME_BITS'd117933461, `RNS_PRIME_BITS'd969770317, `RNS_PRIME_BITS'd910514587, `RNS_PRIME_BITS'd1527045567, `RNS_PRIME_BITS'd995691261, `RNS_PRIME_BITS'd1948577607, `RNS_PRIME_BITS'd2145706332},
			'{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd666736173, `RNS_PRIME_BITS'd1304369445, `RNS_PRIME_BITS'd1794528825, `RNS_PRIME_BITS'd1499159832, `RNS_PRIME_BITS'd1028696567, `RNS_PRIME_BITS'd1450607929, `RNS_PRIME_BITS'd1252106799, `RNS_PRIME_BITS'd1474879344, `RNS_PRIME_BITS'd844595214, `RNS_PRIME_BITS'd1533898817},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd454755607, `RNS_PRIME_BITS'd1796387302, `RNS_PRIME_BITS'd2065247697, `RNS_PRIME_BITS'd1500655679, `RNS_PRIME_BITS'd1220593693, `RNS_PRIME_BITS'd791961431, `RNS_PRIME_BITS'd643624714, `RNS_PRIME_BITS'd488697640, `RNS_PRIME_BITS'd1500839681, `RNS_PRIME_BITS'd924337029},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd1381211600, `RNS_PRIME_BITS'd198408738, `RNS_PRIME_BITS'd469876991, `RNS_PRIME_BITS'd771797900, `RNS_PRIME_BITS'd2023901111, `RNS_PRIME_BITS'd1534964215, `RNS_PRIME_BITS'd1564825573, `RNS_PRIME_BITS'd183705654, `RNS_PRIME_BITS'd766371205, `RNS_PRIME_BITS'd1546765752},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd254707800, `RNS_PRIME_BITS'd469169516, `RNS_PRIME_BITS'd1919147771, `RNS_PRIME_BITS'd211225428, `RNS_PRIME_BITS'd866745833, `RNS_PRIME_BITS'd1755399791, `RNS_PRIME_BITS'd1134167816, `RNS_PRIME_BITS'd783514644, `RNS_PRIME_BITS'd1104096838, `RNS_PRIME_BITS'd738589978},
			'{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd2105365369, `RNS_PRIME_BITS'd410412306, `RNS_PRIME_BITS'd1903206157, `RNS_PRIME_BITS'd907075430, `RNS_PRIME_BITS'd665760695, `RNS_PRIME_BITS'd383524058, `RNS_PRIME_BITS'd2095082691, `RNS_PRIME_BITS'd1089120267, `RNS_PRIME_BITS'd36791421, `RNS_PRIME_BITS'd1689620762},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd816978877, `RNS_PRIME_BITS'd1740930797, `RNS_PRIME_BITS'd388955725, `RNS_PRIME_BITS'd1531118562, `RNS_PRIME_BITS'd1377044326, `RNS_PRIME_BITS'd169254052, `RNS_PRIME_BITS'd907014959, `RNS_PRIME_BITS'd2024070620, `RNS_PRIME_BITS'd2001497750, `RNS_PRIME_BITS'd772430705},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd1337979240, `RNS_PRIME_BITS'd1347938008, `RNS_PRIME_BITS'd22345998, `RNS_PRIME_BITS'd2067964738, `RNS_PRIME_BITS'd1101885111, `RNS_PRIME_BITS'd1334025046, `RNS_PRIME_BITS'd1599461484, `RNS_PRIME_BITS'd217589556, `RNS_PRIME_BITS'd845242412, `RNS_PRIME_BITS'd1115974534},
			'{`RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd1167248610, `RNS_PRIME_BITS'd1603490954, `RNS_PRIME_BITS'd170665898, `RNS_PRIME_BITS'd981588349, `RNS_PRIME_BITS'd469649202, `RNS_PRIME_BITS'd451812643, `RNS_PRIME_BITS'd1073036117, `RNS_PRIME_BITS'd276585797, `RNS_PRIME_BITS'd237334585, `RNS_PRIME_BITS'd2147254786},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd544595951, `RNS_PRIME_BITS'd332844411, `RNS_PRIME_BITS'd2044024803, `RNS_PRIME_BITS'd1017817074, `RNS_PRIME_BITS'd50582275, `RNS_PRIME_BITS'd1274274425, `RNS_PRIME_BITS'd941795823, `RNS_PRIME_BITS'd866674053, `RNS_PRIME_BITS'd1046301558, `RNS_PRIME_BITS'd1482666159},
			'{`RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd1071308433, `RNS_PRIME_BITS'd177120984, `RNS_PRIME_BITS'd1181274533, `RNS_PRIME_BITS'd545498313, `RNS_PRIME_BITS'd1182354334, `RNS_PRIME_BITS'd142722001, `RNS_PRIME_BITS'd1109512168, `RNS_PRIME_BITS'd992164114, `RNS_PRIME_BITS'd1936572605, `RNS_PRIME_BITS'd733223811},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd633297840, `RNS_PRIME_BITS'd1642317120, `RNS_PRIME_BITS'd632356005, `RNS_PRIME_BITS'd287441253, `RNS_PRIME_BITS'd1053162745, `RNS_PRIME_BITS'd849196473, `RNS_PRIME_BITS'd1988190551, `RNS_PRIME_BITS'd1352762144, `RNS_PRIME_BITS'd1936458115, `RNS_PRIME_BITS'd331985327}
		},
		'{
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1071949173, `RNS_PRIME_BITS'd183117999, `RNS_PRIME_BITS'd1887400053, `RNS_PRIME_BITS'd1376158118, `RNS_PRIME_BITS'd1629179269, `RNS_PRIME_BITS'd826092867, `RNS_PRIME_BITS'd1888200167, `RNS_PRIME_BITS'd336173160, `RNS_PRIME_BITS'd21289048, `RNS_PRIME_BITS'd1978400453},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1674372888, `RNS_PRIME_BITS'd446719271, `RNS_PRIME_BITS'd1053760783, `RNS_PRIME_BITS'd1756598555, `RNS_PRIME_BITS'd456433363, `RNS_PRIME_BITS'd923272630, `RNS_PRIME_BITS'd620854330, `RNS_PRIME_BITS'd1409282053, `RNS_PRIME_BITS'd808197817, `RNS_PRIME_BITS'd619006815},
			'{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd1260773675, `RNS_PRIME_BITS'd1580716284, `RNS_PRIME_BITS'd625403534, `RNS_PRIME_BITS'd591266689, `RNS_PRIME_BITS'd1739304459, `RNS_PRIME_BITS'd561545882, `RNS_PRIME_BITS'd7491407, `RNS_PRIME_BITS'd95098928, `RNS_PRIME_BITS'd491026664, `RNS_PRIME_BITS'd606462801},
			'{`RNS_PRIME_BITS'd156, `RNS_PRIME_BITS'd1186602152, `RNS_PRIME_BITS'd1659474382, `RNS_PRIME_BITS'd1569761478, `RNS_PRIME_BITS'd951576757, `RNS_PRIME_BITS'd1836439901, `RNS_PRIME_BITS'd796050041, `RNS_PRIME_BITS'd1463486788, `RNS_PRIME_BITS'd2042018018, `RNS_PRIME_BITS'd1148989093, `RNS_PRIME_BITS'd510666746},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1742169867, `RNS_PRIME_BITS'd1488570758, `RNS_PRIME_BITS'd1900863933, `RNS_PRIME_BITS'd813006813, `RNS_PRIME_BITS'd1186795612, `RNS_PRIME_BITS'd116046918, `RNS_PRIME_BITS'd432469312, `RNS_PRIME_BITS'd1074965162, `RNS_PRIME_BITS'd2090238844, `RNS_PRIME_BITS'd1476590174},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd74359362, `RNS_PRIME_BITS'd116494425, `RNS_PRIME_BITS'd1772450492, `RNS_PRIME_BITS'd2113184363, `RNS_PRIME_BITS'd1731817852, `RNS_PRIME_BITS'd802787944, `RNS_PRIME_BITS'd1141689633, `RNS_PRIME_BITS'd830427413, `RNS_PRIME_BITS'd1249413134, `RNS_PRIME_BITS'd958286481},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd1777387860, `RNS_PRIME_BITS'd1569171508, `RNS_PRIME_BITS'd1441865977, `RNS_PRIME_BITS'd136216553, `RNS_PRIME_BITS'd480776430, `RNS_PRIME_BITS'd2025831634, `RNS_PRIME_BITS'd2013461358, `RNS_PRIME_BITS'd444798078, `RNS_PRIME_BITS'd22203557, `RNS_PRIME_BITS'd110537304},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd1037117329, `RNS_PRIME_BITS'd1429764733, `RNS_PRIME_BITS'd874435822, `RNS_PRIME_BITS'd1874557671, `RNS_PRIME_BITS'd598969008, `RNS_PRIME_BITS'd1763092166, `RNS_PRIME_BITS'd57787589, `RNS_PRIME_BITS'd1318554027, `RNS_PRIME_BITS'd1042421178, `RNS_PRIME_BITS'd2145911719},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd1160577968, `RNS_PRIME_BITS'd794134712, `RNS_PRIME_BITS'd1886024178, `RNS_PRIME_BITS'd809969255, `RNS_PRIME_BITS'd1655258816, `RNS_PRIME_BITS'd1522193282, `RNS_PRIME_BITS'd1924101425, `RNS_PRIME_BITS'd1979068380, `RNS_PRIME_BITS'd1189943286, `RNS_PRIME_BITS'd2129372632},
			'{`RNS_PRIME_BITS'd65, `RNS_PRIME_BITS'd262793099, `RNS_PRIME_BITS'd2121929895, `RNS_PRIME_BITS'd2077486483, `RNS_PRIME_BITS'd1873944392, `RNS_PRIME_BITS'd1206540732, `RNS_PRIME_BITS'd2122399069, `RNS_PRIME_BITS'd1457870051, `RNS_PRIME_BITS'd450697652, `RNS_PRIME_BITS'd832613448, `RNS_PRIME_BITS'd1317130181},
			'{`RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd1346895426, `RNS_PRIME_BITS'd369958396, `RNS_PRIME_BITS'd990162012, `RNS_PRIME_BITS'd1637148926, `RNS_PRIME_BITS'd656083518, `RNS_PRIME_BITS'd1842513321, `RNS_PRIME_BITS'd937941792, `RNS_PRIME_BITS'd2016162590, `RNS_PRIME_BITS'd1513212193, `RNS_PRIME_BITS'd1383102411},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1877975351, `RNS_PRIME_BITS'd116059990, `RNS_PRIME_BITS'd347919052, `RNS_PRIME_BITS'd1261437484, `RNS_PRIME_BITS'd2033607336, `RNS_PRIME_BITS'd961784740, `RNS_PRIME_BITS'd1369784752, `RNS_PRIME_BITS'd156219139, `RNS_PRIME_BITS'd701776419, `RNS_PRIME_BITS'd668674341},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd1694799654, `RNS_PRIME_BITS'd2123545879, `RNS_PRIME_BITS'd1845290585, `RNS_PRIME_BITS'd1808719056, `RNS_PRIME_BITS'd506150510, `RNS_PRIME_BITS'd1630663733, `RNS_PRIME_BITS'd504489429, `RNS_PRIME_BITS'd407956393, `RNS_PRIME_BITS'd578715436, `RNS_PRIME_BITS'd1273276830},
			'{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd256637348, `RNS_PRIME_BITS'd1445529899, `RNS_PRIME_BITS'd935835327, `RNS_PRIME_BITS'd1040375247, `RNS_PRIME_BITS'd179402422, `RNS_PRIME_BITS'd1433937734, `RNS_PRIME_BITS'd1017988555, `RNS_PRIME_BITS'd1179783156, `RNS_PRIME_BITS'd617324358, `RNS_PRIME_BITS'd1830025915},
			'{`RNS_PRIME_BITS'd6, `RNS_PRIME_BITS'd847675295, `RNS_PRIME_BITS'd1339973626, `RNS_PRIME_BITS'd1728772871, `RNS_PRIME_BITS'd620488165, `RNS_PRIME_BITS'd642903007, `RNS_PRIME_BITS'd178009753, `RNS_PRIME_BITS'd224091063, `RNS_PRIME_BITS'd2072622053, `RNS_PRIME_BITS'd1463553277, `RNS_PRIME_BITS'd1922708575},
			'{`RNS_PRIME_BITS'd210, `RNS_PRIME_BITS'd922425555, `RNS_PRIME_BITS'd401772308, `RNS_PRIME_BITS'd960209100, `RNS_PRIME_BITS'd1294905795, `RNS_PRIME_BITS'd743795939, `RNS_PRIME_BITS'd946449119, `RNS_PRIME_BITS'd612106984, `RNS_PRIME_BITS'd795256685, `RNS_PRIME_BITS'd1180296917, `RNS_PRIME_BITS'd1186589394},
			'{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd1428592465, `RNS_PRIME_BITS'd502048311, `RNS_PRIME_BITS'd677059007, `RNS_PRIME_BITS'd1034905853, `RNS_PRIME_BITS'd1537090939, `RNS_PRIME_BITS'd1198179598, `RNS_PRIME_BITS'd1143418979, `RNS_PRIME_BITS'd520493764, `RNS_PRIME_BITS'd1987428434, `RNS_PRIME_BITS'd716823501},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd371156343, `RNS_PRIME_BITS'd1403383334, `RNS_PRIME_BITS'd886194300, `RNS_PRIME_BITS'd1190923666, `RNS_PRIME_BITS'd1206654267, `RNS_PRIME_BITS'd1820900288, `RNS_PRIME_BITS'd1502959195, `RNS_PRIME_BITS'd1977323623, `RNS_PRIME_BITS'd1932445697, `RNS_PRIME_BITS'd1649310753},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd882905420, `RNS_PRIME_BITS'd1864380162, `RNS_PRIME_BITS'd1361363561, `RNS_PRIME_BITS'd56512039, `RNS_PRIME_BITS'd1252720722, `RNS_PRIME_BITS'd206434474, `RNS_PRIME_BITS'd1695276021, `RNS_PRIME_BITS'd1253490274, `RNS_PRIME_BITS'd1402784099, `RNS_PRIME_BITS'd21326092},
			'{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd1709050824, `RNS_PRIME_BITS'd1496333282, `RNS_PRIME_BITS'd669220115, `RNS_PRIME_BITS'd2073935571, `RNS_PRIME_BITS'd1416320280, `RNS_PRIME_BITS'd187286800, `RNS_PRIME_BITS'd7606038, `RNS_PRIME_BITS'd758238598, `RNS_PRIME_BITS'd1532662942, `RNS_PRIME_BITS'd2023175823},
			'{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd1578221698, `RNS_PRIME_BITS'd1677218639, `RNS_PRIME_BITS'd1398064352, `RNS_PRIME_BITS'd1109686688, `RNS_PRIME_BITS'd234920308, `RNS_PRIME_BITS'd660020838, `RNS_PRIME_BITS'd1984551441, `RNS_PRIME_BITS'd2029009578, `RNS_PRIME_BITS'd1810077466, `RNS_PRIME_BITS'd1611309010},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd407223402, `RNS_PRIME_BITS'd1602868668, `RNS_PRIME_BITS'd260865472, `RNS_PRIME_BITS'd1183690885, `RNS_PRIME_BITS'd1522818180, `RNS_PRIME_BITS'd1672347026, `RNS_PRIME_BITS'd1997054979, `RNS_PRIME_BITS'd439377839, `RNS_PRIME_BITS'd1407862169, `RNS_PRIME_BITS'd987820074},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd311363603, `RNS_PRIME_BITS'd454174774, `RNS_PRIME_BITS'd1308547036, `RNS_PRIME_BITS'd101398299, `RNS_PRIME_BITS'd1130712339, `RNS_PRIME_BITS'd1017979193, `RNS_PRIME_BITS'd1659080984, `RNS_PRIME_BITS'd359261879, `RNS_PRIME_BITS'd27527951, `RNS_PRIME_BITS'd1577869248},
			'{`RNS_PRIME_BITS'd169, `RNS_PRIME_BITS'd1994202050, `RNS_PRIME_BITS'd812168176, `RNS_PRIME_BITS'd21870459, `RNS_PRIME_BITS'd2043256972, `RNS_PRIME_BITS'd1039874137, `RNS_PRIME_BITS'd2039083825, `RNS_PRIME_BITS'd964657090, `RNS_PRIME_BITS'd1616679478, `RNS_PRIME_BITS'd1665630174, `RNS_PRIME_BITS'd2091417461},
			'{`RNS_PRIME_BITS'd170, `RNS_PRIME_BITS'd1183765700, `RNS_PRIME_BITS'd1910652704, `RNS_PRIME_BITS'd1132466554, `RNS_PRIME_BITS'd268483656, `RNS_PRIME_BITS'd484338396, `RNS_PRIME_BITS'd512825741, `RNS_PRIME_BITS'd785015160, `RNS_PRIME_BITS'd1529914929, `RNS_PRIME_BITS'd1784855229, `RNS_PRIME_BITS'd757319094},
			'{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd429128011, `RNS_PRIME_BITS'd1387212799, `RNS_PRIME_BITS'd1806682042, `RNS_PRIME_BITS'd1268700113, `RNS_PRIME_BITS'd1324308382, `RNS_PRIME_BITS'd652259610, `RNS_PRIME_BITS'd1418774986, `RNS_PRIME_BITS'd1719028740, `RNS_PRIME_BITS'd2105730329, `RNS_PRIME_BITS'd885930301},
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd638539241, `RNS_PRIME_BITS'd1524040504, `RNS_PRIME_BITS'd465441772, `RNS_PRIME_BITS'd45045752, `RNS_PRIME_BITS'd1087220352, `RNS_PRIME_BITS'd1742785056, `RNS_PRIME_BITS'd1781350150, `RNS_PRIME_BITS'd1481437797, `RNS_PRIME_BITS'd1109010764, `RNS_PRIME_BITS'd1609778726},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd2027168079, `RNS_PRIME_BITS'd1894667374, `RNS_PRIME_BITS'd267234932, `RNS_PRIME_BITS'd1000155678, `RNS_PRIME_BITS'd874343171, `RNS_PRIME_BITS'd461943072, `RNS_PRIME_BITS'd524900293, `RNS_PRIME_BITS'd233096531, `RNS_PRIME_BITS'd1843356303, `RNS_PRIME_BITS'd133288502},
			'{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd2138839197, `RNS_PRIME_BITS'd1958475766, `RNS_PRIME_BITS'd2093896265, `RNS_PRIME_BITS'd1043136997, `RNS_PRIME_BITS'd1615286639, `RNS_PRIME_BITS'd1130676792, `RNS_PRIME_BITS'd1706004929, `RNS_PRIME_BITS'd1503498928, `RNS_PRIME_BITS'd191968825, `RNS_PRIME_BITS'd1056633049},
			'{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd789307144, `RNS_PRIME_BITS'd823163169, `RNS_PRIME_BITS'd717872639, `RNS_PRIME_BITS'd557776342, `RNS_PRIME_BITS'd1308477027, `RNS_PRIME_BITS'd1969268214, `RNS_PRIME_BITS'd362237114, `RNS_PRIME_BITS'd2049542735, `RNS_PRIME_BITS'd100563678, `RNS_PRIME_BITS'd422786923},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd2037555191, `RNS_PRIME_BITS'd928036423, `RNS_PRIME_BITS'd2022884891, `RNS_PRIME_BITS'd1599851167, `RNS_PRIME_BITS'd1281229743, `RNS_PRIME_BITS'd1067017411, `RNS_PRIME_BITS'd1695836816, `RNS_PRIME_BITS'd82471313, `RNS_PRIME_BITS'd1399392295, `RNS_PRIME_BITS'd424188337},
			'{`RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd1488753794, `RNS_PRIME_BITS'd304910566, `RNS_PRIME_BITS'd1710234530, `RNS_PRIME_BITS'd883824648, `RNS_PRIME_BITS'd1785889672, `RNS_PRIME_BITS'd1569111768, `RNS_PRIME_BITS'd304037453, `RNS_PRIME_BITS'd1755635575, `RNS_PRIME_BITS'd1811147510, `RNS_PRIME_BITS'd2019360265},
			'{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd1134831169, `RNS_PRIME_BITS'd1467998358, `RNS_PRIME_BITS'd715727843, `RNS_PRIME_BITS'd1081079509, `RNS_PRIME_BITS'd182350517, `RNS_PRIME_BITS'd1634912862, `RNS_PRIME_BITS'd1898535294, `RNS_PRIME_BITS'd760571975, `RNS_PRIME_BITS'd567268552, `RNS_PRIME_BITS'd128751838},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd2112122460, `RNS_PRIME_BITS'd8113561, `RNS_PRIME_BITS'd1978367443, `RNS_PRIME_BITS'd885878873, `RNS_PRIME_BITS'd1054154075, `RNS_PRIME_BITS'd734701926, `RNS_PRIME_BITS'd778830896, `RNS_PRIME_BITS'd614686835, `RNS_PRIME_BITS'd903107778, `RNS_PRIME_BITS'd167770899},
			'{`RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd225279763, `RNS_PRIME_BITS'd329267680, `RNS_PRIME_BITS'd869433125, `RNS_PRIME_BITS'd92649644, `RNS_PRIME_BITS'd1956902978, `RNS_PRIME_BITS'd335341295, `RNS_PRIME_BITS'd95732843, `RNS_PRIME_BITS'd1888439119, `RNS_PRIME_BITS'd856834203, `RNS_PRIME_BITS'd1270498048},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1035876073, `RNS_PRIME_BITS'd593618531, `RNS_PRIME_BITS'd119278412, `RNS_PRIME_BITS'd425887380, `RNS_PRIME_BITS'd57859843, `RNS_PRIME_BITS'd430428972, `RNS_PRIME_BITS'd1110930763, `RNS_PRIME_BITS'd1937258344, `RNS_PRIME_BITS'd388394255, `RNS_PRIME_BITS'd60585110},
			'{`RNS_PRIME_BITS'd190, `RNS_PRIME_BITS'd314198983, `RNS_PRIME_BITS'd1784689567, `RNS_PRIME_BITS'd1078242304, `RNS_PRIME_BITS'd1770708593, `RNS_PRIME_BITS'd1238202625, `RNS_PRIME_BITS'd2071219325, `RNS_PRIME_BITS'd376170328, `RNS_PRIME_BITS'd1221608071, `RNS_PRIME_BITS'd99779297, `RNS_PRIME_BITS'd1500123181},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1922925644, `RNS_PRIME_BITS'd1440861228, `RNS_PRIME_BITS'd315941632, `RNS_PRIME_BITS'd1537420147, `RNS_PRIME_BITS'd1387578946, `RNS_PRIME_BITS'd388271832, `RNS_PRIME_BITS'd920614593, `RNS_PRIME_BITS'd1192636634, `RNS_PRIME_BITS'd582903, `RNS_PRIME_BITS'd25516772},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd514100804, `RNS_PRIME_BITS'd1319147413, `RNS_PRIME_BITS'd1152001911, `RNS_PRIME_BITS'd298842349, `RNS_PRIME_BITS'd1656248434, `RNS_PRIME_BITS'd1246074280, `RNS_PRIME_BITS'd1811833943, `RNS_PRIME_BITS'd580732723, `RNS_PRIME_BITS'd1883342472, `RNS_PRIME_BITS'd1534416785},
			'{`RNS_PRIME_BITS'd32, `RNS_PRIME_BITS'd205344120, `RNS_PRIME_BITS'd585840830, `RNS_PRIME_BITS'd1180576594, `RNS_PRIME_BITS'd115398121, `RNS_PRIME_BITS'd1014965676, `RNS_PRIME_BITS'd486202073, `RNS_PRIME_BITS'd904561231, `RNS_PRIME_BITS'd1040642742, `RNS_PRIME_BITS'd292627552, `RNS_PRIME_BITS'd1636738649},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd1674258249, `RNS_PRIME_BITS'd1494623564, `RNS_PRIME_BITS'd1687956038, `RNS_PRIME_BITS'd1503345269, `RNS_PRIME_BITS'd1237948697, `RNS_PRIME_BITS'd1904398235, `RNS_PRIME_BITS'd744383252, `RNS_PRIME_BITS'd114004353, `RNS_PRIME_BITS'd1934553852, `RNS_PRIME_BITS'd965879722},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd686425061, `RNS_PRIME_BITS'd709618911, `RNS_PRIME_BITS'd257366225, `RNS_PRIME_BITS'd559133558, `RNS_PRIME_BITS'd972588978, `RNS_PRIME_BITS'd1723588688, `RNS_PRIME_BITS'd1900587433, `RNS_PRIME_BITS'd392119190, `RNS_PRIME_BITS'd170746619, `RNS_PRIME_BITS'd1942963090},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd318359049, `RNS_PRIME_BITS'd1664680159, `RNS_PRIME_BITS'd664204501, `RNS_PRIME_BITS'd1919608803, `RNS_PRIME_BITS'd843079740, `RNS_PRIME_BITS'd610865944, `RNS_PRIME_BITS'd209551215, `RNS_PRIME_BITS'd438475805, `RNS_PRIME_BITS'd278984482, `RNS_PRIME_BITS'd1674350665},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd1360647303, `RNS_PRIME_BITS'd1708701190, `RNS_PRIME_BITS'd1210454273, `RNS_PRIME_BITS'd1832054185, `RNS_PRIME_BITS'd1052903264, `RNS_PRIME_BITS'd128077122, `RNS_PRIME_BITS'd975280264, `RNS_PRIME_BITS'd1267912710, `RNS_PRIME_BITS'd746763716, `RNS_PRIME_BITS'd1764420488},
			'{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd961202458, `RNS_PRIME_BITS'd789436046, `RNS_PRIME_BITS'd1532553559, `RNS_PRIME_BITS'd557337327, `RNS_PRIME_BITS'd1702447767, `RNS_PRIME_BITS'd1869387258, `RNS_PRIME_BITS'd991781017, `RNS_PRIME_BITS'd599971478, `RNS_PRIME_BITS'd1984485596, `RNS_PRIME_BITS'd1229967891},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd1680380819, `RNS_PRIME_BITS'd490617682, `RNS_PRIME_BITS'd134909027, `RNS_PRIME_BITS'd1454993387, `RNS_PRIME_BITS'd1463760555, `RNS_PRIME_BITS'd176472365, `RNS_PRIME_BITS'd405165357, `RNS_PRIME_BITS'd1909250531, `RNS_PRIME_BITS'd463892239, `RNS_PRIME_BITS'd1962383673},
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd2065249957, `RNS_PRIME_BITS'd1076970720, `RNS_PRIME_BITS'd1745332931, `RNS_PRIME_BITS'd165790248, `RNS_PRIME_BITS'd122040332, `RNS_PRIME_BITS'd1537145013, `RNS_PRIME_BITS'd336868885, `RNS_PRIME_BITS'd431877522, `RNS_PRIME_BITS'd733175249, `RNS_PRIME_BITS'd898591109},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd743436892, `RNS_PRIME_BITS'd304757575, `RNS_PRIME_BITS'd2070374395, `RNS_PRIME_BITS'd1887651520, `RNS_PRIME_BITS'd2017164177, `RNS_PRIME_BITS'd2139440781, `RNS_PRIME_BITS'd1453004132, `RNS_PRIME_BITS'd464668391, `RNS_PRIME_BITS'd1885318016, `RNS_PRIME_BITS'd1518882868},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd2122524636, `RNS_PRIME_BITS'd529106586, `RNS_PRIME_BITS'd739559141, `RNS_PRIME_BITS'd1435958920, `RNS_PRIME_BITS'd823906974, `RNS_PRIME_BITS'd1781996288, `RNS_PRIME_BITS'd1683077951, `RNS_PRIME_BITS'd2007352462, `RNS_PRIME_BITS'd259587288, `RNS_PRIME_BITS'd334830297},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd899556659, `RNS_PRIME_BITS'd202300419, `RNS_PRIME_BITS'd220099240, `RNS_PRIME_BITS'd446504188, `RNS_PRIME_BITS'd2067954051, `RNS_PRIME_BITS'd1913247950, `RNS_PRIME_BITS'd1518924337, `RNS_PRIME_BITS'd51763429, `RNS_PRIME_BITS'd995086604, `RNS_PRIME_BITS'd2006765849},
			'{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd2027638776, `RNS_PRIME_BITS'd1244077455, `RNS_PRIME_BITS'd479941227, `RNS_PRIME_BITS'd110902033, `RNS_PRIME_BITS'd862373901, `RNS_PRIME_BITS'd1362451662, `RNS_PRIME_BITS'd1540325228, `RNS_PRIME_BITS'd2028138797, `RNS_PRIME_BITS'd558858150, `RNS_PRIME_BITS'd519845124},
			'{`RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd407698325, `RNS_PRIME_BITS'd1363931285, `RNS_PRIME_BITS'd1198127103, `RNS_PRIME_BITS'd115262392, `RNS_PRIME_BITS'd1163827239, `RNS_PRIME_BITS'd114862328, `RNS_PRIME_BITS'd848117678, `RNS_PRIME_BITS'd707647524, `RNS_PRIME_BITS'd447704888, `RNS_PRIME_BITS'd1803961406},
			'{`RNS_PRIME_BITS'd125, `RNS_PRIME_BITS'd770222703, `RNS_PRIME_BITS'd538184517, `RNS_PRIME_BITS'd775897995, `RNS_PRIME_BITS'd1470802220, `RNS_PRIME_BITS'd2056478144, `RNS_PRIME_BITS'd1950551324, `RNS_PRIME_BITS'd288293387, `RNS_PRIME_BITS'd798964000, `RNS_PRIME_BITS'd788795025, `RNS_PRIME_BITS'd1847860586},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd753228863, `RNS_PRIME_BITS'd1240611315, `RNS_PRIME_BITS'd550916918, `RNS_PRIME_BITS'd734119173, `RNS_PRIME_BITS'd554674391, `RNS_PRIME_BITS'd260850260, `RNS_PRIME_BITS'd2027835604, `RNS_PRIME_BITS'd2076154964, `RNS_PRIME_BITS'd1815281712, `RNS_PRIME_BITS'd377262698},
			'{`RNS_PRIME_BITS'd22, `RNS_PRIME_BITS'd1677321334, `RNS_PRIME_BITS'd800774920, `RNS_PRIME_BITS'd1851656598, `RNS_PRIME_BITS'd416528655, `RNS_PRIME_BITS'd999449317, `RNS_PRIME_BITS'd1590323900, `RNS_PRIME_BITS'd1142943505, `RNS_PRIME_BITS'd149267225, `RNS_PRIME_BITS'd1064893194, `RNS_PRIME_BITS'd1239088933},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd417014783, `RNS_PRIME_BITS'd1971564584, `RNS_PRIME_BITS'd1346005350, `RNS_PRIME_BITS'd1791908716, `RNS_PRIME_BITS'd76427620, `RNS_PRIME_BITS'd1284013218, `RNS_PRIME_BITS'd2098565772, `RNS_PRIME_BITS'd1446565664, `RNS_PRIME_BITS'd1163270812, `RNS_PRIME_BITS'd1640747149},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd1580559365, `RNS_PRIME_BITS'd719037426, `RNS_PRIME_BITS'd275571075, `RNS_PRIME_BITS'd930128443, `RNS_PRIME_BITS'd1091007418, `RNS_PRIME_BITS'd970824606, `RNS_PRIME_BITS'd40954432, `RNS_PRIME_BITS'd1781855541, `RNS_PRIME_BITS'd951124184, `RNS_PRIME_BITS'd1321331437},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd1107680624, `RNS_PRIME_BITS'd995884756, `RNS_PRIME_BITS'd284183636, `RNS_PRIME_BITS'd1995089114, `RNS_PRIME_BITS'd1672315130, `RNS_PRIME_BITS'd1924781693, `RNS_PRIME_BITS'd878115010, `RNS_PRIME_BITS'd259794964, `RNS_PRIME_BITS'd834287783, `RNS_PRIME_BITS'd893210332},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1186242609, `RNS_PRIME_BITS'd1364729528, `RNS_PRIME_BITS'd40315126, `RNS_PRIME_BITS'd1753211630, `RNS_PRIME_BITS'd813915482, `RNS_PRIME_BITS'd98264556, `RNS_PRIME_BITS'd367427412, `RNS_PRIME_BITS'd257153778, `RNS_PRIME_BITS'd1214957078, `RNS_PRIME_BITS'd1507150523},
			'{`RNS_PRIME_BITS'd210, `RNS_PRIME_BITS'd1404455804, `RNS_PRIME_BITS'd1539592576, `RNS_PRIME_BITS'd1804406358, `RNS_PRIME_BITS'd1189433942, `RNS_PRIME_BITS'd200655382, `RNS_PRIME_BITS'd447031920, `RNS_PRIME_BITS'd495508209, `RNS_PRIME_BITS'd1640572009, `RNS_PRIME_BITS'd683687045, `RNS_PRIME_BITS'd1198265148},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd815611521, `RNS_PRIME_BITS'd222639021, `RNS_PRIME_BITS'd1437067345, `RNS_PRIME_BITS'd1388010570, `RNS_PRIME_BITS'd530241525, `RNS_PRIME_BITS'd1651178178, `RNS_PRIME_BITS'd448856107, `RNS_PRIME_BITS'd1626401454, `RNS_PRIME_BITS'd1252161744, `RNS_PRIME_BITS'd1714893946},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1803691360, `RNS_PRIME_BITS'd2072279921, `RNS_PRIME_BITS'd1037480712, `RNS_PRIME_BITS'd1352233960, `RNS_PRIME_BITS'd1175806607, `RNS_PRIME_BITS'd395898123, `RNS_PRIME_BITS'd1118263484, `RNS_PRIME_BITS'd1795875378, `RNS_PRIME_BITS'd1069520845, `RNS_PRIME_BITS'd204807639},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd2034356509, `RNS_PRIME_BITS'd168983359, `RNS_PRIME_BITS'd1875319407, `RNS_PRIME_BITS'd1900502433, `RNS_PRIME_BITS'd1158503763, `RNS_PRIME_BITS'd379598526, `RNS_PRIME_BITS'd66318495, `RNS_PRIME_BITS'd76535735, `RNS_PRIME_BITS'd1960146339, `RNS_PRIME_BITS'd1199375967},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1396745173, `RNS_PRIME_BITS'd208752612, `RNS_PRIME_BITS'd1576358889, `RNS_PRIME_BITS'd135424037, `RNS_PRIME_BITS'd1110504270, `RNS_PRIME_BITS'd1386083419, `RNS_PRIME_BITS'd865521619, `RNS_PRIME_BITS'd825303066, `RNS_PRIME_BITS'd1807986135, `RNS_PRIME_BITS'd1097834131}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd2120820943, `RNS_PRIME_BITS'd1993896682, `RNS_PRIME_BITS'd504129854, `RNS_PRIME_BITS'd1935907347, `RNS_PRIME_BITS'd1117170337, `RNS_PRIME_BITS'd524162989, `RNS_PRIME_BITS'd1996449838, `RNS_PRIME_BITS'd1523748127, `RNS_PRIME_BITS'd2116676240, `RNS_PRIME_BITS'd951672547},
			'{`RNS_PRIME_BITS'd190, `RNS_PRIME_BITS'd598009359, `RNS_PRIME_BITS'd1050569549, `RNS_PRIME_BITS'd267146485, `RNS_PRIME_BITS'd671323730, `RNS_PRIME_BITS'd1222008356, `RNS_PRIME_BITS'd226786407, `RNS_PRIME_BITS'd809332597, `RNS_PRIME_BITS'd1421607399, `RNS_PRIME_BITS'd1809088231, `RNS_PRIME_BITS'd1267564003},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd733343979, `RNS_PRIME_BITS'd1386461334, `RNS_PRIME_BITS'd244876494, `RNS_PRIME_BITS'd638577846, `RNS_PRIME_BITS'd1807154147, `RNS_PRIME_BITS'd1491848368, `RNS_PRIME_BITS'd1707044273, `RNS_PRIME_BITS'd1339656238, `RNS_PRIME_BITS'd1970449665, `RNS_PRIME_BITS'd921603474},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1800321465, `RNS_PRIME_BITS'd555524051, `RNS_PRIME_BITS'd473991296, `RNS_PRIME_BITS'd341948731, `RNS_PRIME_BITS'd2127994793, `RNS_PRIME_BITS'd1475761216, `RNS_PRIME_BITS'd637343389, `RNS_PRIME_BITS'd411479394, `RNS_PRIME_BITS'd1068739877, `RNS_PRIME_BITS'd2001790556},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd920883317, `RNS_PRIME_BITS'd2075623301, `RNS_PRIME_BITS'd845584306, `RNS_PRIME_BITS'd1532525047, `RNS_PRIME_BITS'd983568479, `RNS_PRIME_BITS'd104272907, `RNS_PRIME_BITS'd1510950855, `RNS_PRIME_BITS'd1391291706, `RNS_PRIME_BITS'd336733398, `RNS_PRIME_BITS'd116814755},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd235233920, `RNS_PRIME_BITS'd551023015, `RNS_PRIME_BITS'd1327026559, `RNS_PRIME_BITS'd1090450089, `RNS_PRIME_BITS'd2134543417, `RNS_PRIME_BITS'd1360184500, `RNS_PRIME_BITS'd1001707131, `RNS_PRIME_BITS'd1578633503, `RNS_PRIME_BITS'd809912994, `RNS_PRIME_BITS'd1422963867},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd125250816, `RNS_PRIME_BITS'd219755185, `RNS_PRIME_BITS'd1471752856, `RNS_PRIME_BITS'd360704811, `RNS_PRIME_BITS'd1164889660, `RNS_PRIME_BITS'd618442700, `RNS_PRIME_BITS'd1578233941, `RNS_PRIME_BITS'd1550555452, `RNS_PRIME_BITS'd1411646224, `RNS_PRIME_BITS'd183402407},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd727012638, `RNS_PRIME_BITS'd1550340675, `RNS_PRIME_BITS'd370097028, `RNS_PRIME_BITS'd1303090563, `RNS_PRIME_BITS'd1548231734, `RNS_PRIME_BITS'd1815733696, `RNS_PRIME_BITS'd529605270, `RNS_PRIME_BITS'd2087391567, `RNS_PRIME_BITS'd376656255, `RNS_PRIME_BITS'd1195726978},
			'{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd361636896, `RNS_PRIME_BITS'd75570555, `RNS_PRIME_BITS'd95407925, `RNS_PRIME_BITS'd540596697, `RNS_PRIME_BITS'd1941684858, `RNS_PRIME_BITS'd889229760, `RNS_PRIME_BITS'd141367125, `RNS_PRIME_BITS'd653628439, `RNS_PRIME_BITS'd1014020786, `RNS_PRIME_BITS'd901127334},
			'{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd745382493, `RNS_PRIME_BITS'd990040693, `RNS_PRIME_BITS'd1582435379, `RNS_PRIME_BITS'd866267702, `RNS_PRIME_BITS'd2097859982, `RNS_PRIME_BITS'd1873305046, `RNS_PRIME_BITS'd1207241132, `RNS_PRIME_BITS'd1274097205, `RNS_PRIME_BITS'd1459662681, `RNS_PRIME_BITS'd232074785},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd34967681, `RNS_PRIME_BITS'd763981419, `RNS_PRIME_BITS'd401623355, `RNS_PRIME_BITS'd797471654, `RNS_PRIME_BITS'd1809331665, `RNS_PRIME_BITS'd719918297, `RNS_PRIME_BITS'd538237392, `RNS_PRIME_BITS'd1874533145, `RNS_PRIME_BITS'd1563210145, `RNS_PRIME_BITS'd202307490},
			'{`RNS_PRIME_BITS'd244, `RNS_PRIME_BITS'd939270925, `RNS_PRIME_BITS'd1512140705, `RNS_PRIME_BITS'd10915210, `RNS_PRIME_BITS'd1244287886, `RNS_PRIME_BITS'd1633879213, `RNS_PRIME_BITS'd178297214, `RNS_PRIME_BITS'd357108422, `RNS_PRIME_BITS'd1566147826, `RNS_PRIME_BITS'd1464705153, `RNS_PRIME_BITS'd1132545440},
			'{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd1390612485, `RNS_PRIME_BITS'd1302177306, `RNS_PRIME_BITS'd1758121190, `RNS_PRIME_BITS'd1040819011, `RNS_PRIME_BITS'd1907125566, `RNS_PRIME_BITS'd221808555, `RNS_PRIME_BITS'd1426095274, `RNS_PRIME_BITS'd1032897949, `RNS_PRIME_BITS'd474400947, `RNS_PRIME_BITS'd1587818295},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd855210237, `RNS_PRIME_BITS'd1827148933, `RNS_PRIME_BITS'd393230333, `RNS_PRIME_BITS'd1646303305, `RNS_PRIME_BITS'd1542853326, `RNS_PRIME_BITS'd1032565750, `RNS_PRIME_BITS'd1522111084, `RNS_PRIME_BITS'd588991151, `RNS_PRIME_BITS'd654233295, `RNS_PRIME_BITS'd1473014984},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd551513978, `RNS_PRIME_BITS'd1981367168, `RNS_PRIME_BITS'd1317736702, `RNS_PRIME_BITS'd354871793, `RNS_PRIME_BITS'd2005046248, `RNS_PRIME_BITS'd264392086, `RNS_PRIME_BITS'd1134675646, `RNS_PRIME_BITS'd185876217, `RNS_PRIME_BITS'd338206625, `RNS_PRIME_BITS'd642731979},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1600502492, `RNS_PRIME_BITS'd1901958531, `RNS_PRIME_BITS'd1840436703, `RNS_PRIME_BITS'd1118505932, `RNS_PRIME_BITS'd1362144635, `RNS_PRIME_BITS'd917432780, `RNS_PRIME_BITS'd218835629, `RNS_PRIME_BITS'd1938486926, `RNS_PRIME_BITS'd1821470653, `RNS_PRIME_BITS'd1939533329},
			'{`RNS_PRIME_BITS'd172, `RNS_PRIME_BITS'd611925890, `RNS_PRIME_BITS'd598805595, `RNS_PRIME_BITS'd245147245, `RNS_PRIME_BITS'd445051514, `RNS_PRIME_BITS'd432005486, `RNS_PRIME_BITS'd978591903, `RNS_PRIME_BITS'd1378460355, `RNS_PRIME_BITS'd682502495, `RNS_PRIME_BITS'd1212020528, `RNS_PRIME_BITS'd312113928},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd2031692872, `RNS_PRIME_BITS'd1211721979, `RNS_PRIME_BITS'd1844776295, `RNS_PRIME_BITS'd181491356, `RNS_PRIME_BITS'd727345772, `RNS_PRIME_BITS'd936003995, `RNS_PRIME_BITS'd395019672, `RNS_PRIME_BITS'd1122931284, `RNS_PRIME_BITS'd556751601, `RNS_PRIME_BITS'd814562036},
			'{`RNS_PRIME_BITS'd56, `RNS_PRIME_BITS'd1069070354, `RNS_PRIME_BITS'd52917659, `RNS_PRIME_BITS'd2110150647, `RNS_PRIME_BITS'd1560785048, `RNS_PRIME_BITS'd73487444, `RNS_PRIME_BITS'd289562615, `RNS_PRIME_BITS'd1664558228, `RNS_PRIME_BITS'd278902020, `RNS_PRIME_BITS'd1480784826, `RNS_PRIME_BITS'd281570321},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1354925414, `RNS_PRIME_BITS'd2016418111, `RNS_PRIME_BITS'd732724944, `RNS_PRIME_BITS'd211187966, `RNS_PRIME_BITS'd114736206, `RNS_PRIME_BITS'd52345819, `RNS_PRIME_BITS'd1432788676, `RNS_PRIME_BITS'd1616873673, `RNS_PRIME_BITS'd1082688111, `RNS_PRIME_BITS'd978760308},
			'{`RNS_PRIME_BITS'd174, `RNS_PRIME_BITS'd1403005974, `RNS_PRIME_BITS'd601354394, `RNS_PRIME_BITS'd2092439469, `RNS_PRIME_BITS'd1709081016, `RNS_PRIME_BITS'd2044905327, `RNS_PRIME_BITS'd1174721429, `RNS_PRIME_BITS'd1808238613, `RNS_PRIME_BITS'd1851869055, `RNS_PRIME_BITS'd516641912, `RNS_PRIME_BITS'd908988667},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd1770307085, `RNS_PRIME_BITS'd1293835144, `RNS_PRIME_BITS'd2142709247, `RNS_PRIME_BITS'd664457449, `RNS_PRIME_BITS'd1797919046, `RNS_PRIME_BITS'd1187630817, `RNS_PRIME_BITS'd315723906, `RNS_PRIME_BITS'd1701791519, `RNS_PRIME_BITS'd732358514, `RNS_PRIME_BITS'd1637729637},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd207371589, `RNS_PRIME_BITS'd1637854372, `RNS_PRIME_BITS'd960024629, `RNS_PRIME_BITS'd1005880048, `RNS_PRIME_BITS'd1166918319, `RNS_PRIME_BITS'd1607497650, `RNS_PRIME_BITS'd1187888368, `RNS_PRIME_BITS'd1178439087, `RNS_PRIME_BITS'd343339332, `RNS_PRIME_BITS'd317499072},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd175679099, `RNS_PRIME_BITS'd1385373733, `RNS_PRIME_BITS'd1630077147, `RNS_PRIME_BITS'd119211155, `RNS_PRIME_BITS'd677818573, `RNS_PRIME_BITS'd1711927275, `RNS_PRIME_BITS'd959244981, `RNS_PRIME_BITS'd2051947895, `RNS_PRIME_BITS'd511563023, `RNS_PRIME_BITS'd908859375},
			'{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd770153874, `RNS_PRIME_BITS'd871240713, `RNS_PRIME_BITS'd1741954427, `RNS_PRIME_BITS'd336684484, `RNS_PRIME_BITS'd355358588, `RNS_PRIME_BITS'd779914681, `RNS_PRIME_BITS'd1395006618, `RNS_PRIME_BITS'd1458265694, `RNS_PRIME_BITS'd559787320, `RNS_PRIME_BITS'd1514508921},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd2089012429, `RNS_PRIME_BITS'd959445134, `RNS_PRIME_BITS'd177588231, `RNS_PRIME_BITS'd468715906, `RNS_PRIME_BITS'd2057018237, `RNS_PRIME_BITS'd1892456125, `RNS_PRIME_BITS'd170267640, `RNS_PRIME_BITS'd1601353119, `RNS_PRIME_BITS'd1797753382, `RNS_PRIME_BITS'd1270919401},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1795496966, `RNS_PRIME_BITS'd1469964673, `RNS_PRIME_BITS'd1080976901, `RNS_PRIME_BITS'd1259915367, `RNS_PRIME_BITS'd303997573, `RNS_PRIME_BITS'd1810659263, `RNS_PRIME_BITS'd825663517, `RNS_PRIME_BITS'd1192068570, `RNS_PRIME_BITS'd298919414, `RNS_PRIME_BITS'd1226592659},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd1889613997, `RNS_PRIME_BITS'd1726612885, `RNS_PRIME_BITS'd1266919353, `RNS_PRIME_BITS'd1740055755, `RNS_PRIME_BITS'd1589994983, `RNS_PRIME_BITS'd1018761043, `RNS_PRIME_BITS'd1649526891, `RNS_PRIME_BITS'd2013409397, `RNS_PRIME_BITS'd1524745814, `RNS_PRIME_BITS'd252055530},
			'{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd1543253018, `RNS_PRIME_BITS'd636688529, `RNS_PRIME_BITS'd699017913, `RNS_PRIME_BITS'd367107799, `RNS_PRIME_BITS'd496466231, `RNS_PRIME_BITS'd578211471, `RNS_PRIME_BITS'd1033342498, `RNS_PRIME_BITS'd16760824, `RNS_PRIME_BITS'd1778838788, `RNS_PRIME_BITS'd65766136},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd62526508, `RNS_PRIME_BITS'd1348350841, `RNS_PRIME_BITS'd337808360, `RNS_PRIME_BITS'd2057951847, `RNS_PRIME_BITS'd1374694162, `RNS_PRIME_BITS'd866464422, `RNS_PRIME_BITS'd166804404, `RNS_PRIME_BITS'd415001160, `RNS_PRIME_BITS'd1444657410, `RNS_PRIME_BITS'd277210931},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd504932930, `RNS_PRIME_BITS'd1968152411, `RNS_PRIME_BITS'd1487228238, `RNS_PRIME_BITS'd2097828867, `RNS_PRIME_BITS'd1042563290, `RNS_PRIME_BITS'd1263146259, `RNS_PRIME_BITS'd1759744203, `RNS_PRIME_BITS'd2036359424, `RNS_PRIME_BITS'd1850747003, `RNS_PRIME_BITS'd1075264979},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd88993638, `RNS_PRIME_BITS'd1488140504, `RNS_PRIME_BITS'd334137996, `RNS_PRIME_BITS'd2023734025, `RNS_PRIME_BITS'd128589050, `RNS_PRIME_BITS'd1871689909, `RNS_PRIME_BITS'd1758385859, `RNS_PRIME_BITS'd76086652, `RNS_PRIME_BITS'd1259787844, `RNS_PRIME_BITS'd506978106},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1071214495, `RNS_PRIME_BITS'd2129331330, `RNS_PRIME_BITS'd1408399510, `RNS_PRIME_BITS'd1050883280, `RNS_PRIME_BITS'd1004954305, `RNS_PRIME_BITS'd982907170, `RNS_PRIME_BITS'd1327388749, `RNS_PRIME_BITS'd12796089, `RNS_PRIME_BITS'd1462281931, `RNS_PRIME_BITS'd716310410},
			'{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd44725851, `RNS_PRIME_BITS'd1359161033, `RNS_PRIME_BITS'd1706536184, `RNS_PRIME_BITS'd1429274330, `RNS_PRIME_BITS'd854378619, `RNS_PRIME_BITS'd1063204935, `RNS_PRIME_BITS'd1038887997, `RNS_PRIME_BITS'd922883037, `RNS_PRIME_BITS'd1524650002, `RNS_PRIME_BITS'd952402643},
			'{`RNS_PRIME_BITS'd238, `RNS_PRIME_BITS'd393289651, `RNS_PRIME_BITS'd1796417573, `RNS_PRIME_BITS'd819423349, `RNS_PRIME_BITS'd166034118, `RNS_PRIME_BITS'd1605422017, `RNS_PRIME_BITS'd1767495533, `RNS_PRIME_BITS'd2117970759, `RNS_PRIME_BITS'd206637107, `RNS_PRIME_BITS'd376272369, `RNS_PRIME_BITS'd868082014},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1270536485, `RNS_PRIME_BITS'd1191300387, `RNS_PRIME_BITS'd186588943, `RNS_PRIME_BITS'd1807495168, `RNS_PRIME_BITS'd1223577142, `RNS_PRIME_BITS'd563996102, `RNS_PRIME_BITS'd1639794050, `RNS_PRIME_BITS'd1486996066, `RNS_PRIME_BITS'd291661409, `RNS_PRIME_BITS'd1192282578},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1891350802, `RNS_PRIME_BITS'd294607952, `RNS_PRIME_BITS'd954639017, `RNS_PRIME_BITS'd499751311, `RNS_PRIME_BITS'd1019122261, `RNS_PRIME_BITS'd1991399075, `RNS_PRIME_BITS'd1515551961, `RNS_PRIME_BITS'd1600329128, `RNS_PRIME_BITS'd2139923631, `RNS_PRIME_BITS'd145023483},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd973394208, `RNS_PRIME_BITS'd1934502260, `RNS_PRIME_BITS'd65407986, `RNS_PRIME_BITS'd1036591722, `RNS_PRIME_BITS'd312333938, `RNS_PRIME_BITS'd314813529, `RNS_PRIME_BITS'd1512690457, `RNS_PRIME_BITS'd1393037682, `RNS_PRIME_BITS'd1668397107, `RNS_PRIME_BITS'd1040797251},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd882841059, `RNS_PRIME_BITS'd221134310, `RNS_PRIME_BITS'd1528573790, `RNS_PRIME_BITS'd1166485638, `RNS_PRIME_BITS'd1520070977, `RNS_PRIME_BITS'd1344111873, `RNS_PRIME_BITS'd195028482, `RNS_PRIME_BITS'd1164325477, `RNS_PRIME_BITS'd1897879746, `RNS_PRIME_BITS'd1521619094},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd1394052831, `RNS_PRIME_BITS'd1195074954, `RNS_PRIME_BITS'd57757373, `RNS_PRIME_BITS'd1984294396, `RNS_PRIME_BITS'd460968696, `RNS_PRIME_BITS'd1808198494, `RNS_PRIME_BITS'd2072677552, `RNS_PRIME_BITS'd990336370, `RNS_PRIME_BITS'd1494050264, `RNS_PRIME_BITS'd1638989864},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1465514874, `RNS_PRIME_BITS'd445758225, `RNS_PRIME_BITS'd411068779, `RNS_PRIME_BITS'd2121610123, `RNS_PRIME_BITS'd1691831647, `RNS_PRIME_BITS'd2043973417, `RNS_PRIME_BITS'd1724875196, `RNS_PRIME_BITS'd737485154, `RNS_PRIME_BITS'd1811908764, `RNS_PRIME_BITS'd54896738},
			'{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd587317000, `RNS_PRIME_BITS'd1533474935, `RNS_PRIME_BITS'd1788218947, `RNS_PRIME_BITS'd1525661166, `RNS_PRIME_BITS'd801760402, `RNS_PRIME_BITS'd349715315, `RNS_PRIME_BITS'd1816995443, `RNS_PRIME_BITS'd318797850, `RNS_PRIME_BITS'd1375542911, `RNS_PRIME_BITS'd747267757},
			'{`RNS_PRIME_BITS'd204, `RNS_PRIME_BITS'd1854969759, `RNS_PRIME_BITS'd371040217, `RNS_PRIME_BITS'd5208759, `RNS_PRIME_BITS'd690251722, `RNS_PRIME_BITS'd97570762, `RNS_PRIME_BITS'd144573289, `RNS_PRIME_BITS'd553941538, `RNS_PRIME_BITS'd1492013063, `RNS_PRIME_BITS'd1205644364, `RNS_PRIME_BITS'd1731430292},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1928815036, `RNS_PRIME_BITS'd835181530, `RNS_PRIME_BITS'd2001011205, `RNS_PRIME_BITS'd231578252, `RNS_PRIME_BITS'd929967474, `RNS_PRIME_BITS'd210223841, `RNS_PRIME_BITS'd1975714944, `RNS_PRIME_BITS'd394507806, `RNS_PRIME_BITS'd354972718, `RNS_PRIME_BITS'd296985379},
			'{`RNS_PRIME_BITS'd105, `RNS_PRIME_BITS'd1487719583, `RNS_PRIME_BITS'd496160028, `RNS_PRIME_BITS'd981699760, `RNS_PRIME_BITS'd1919706628, `RNS_PRIME_BITS'd1614994336, `RNS_PRIME_BITS'd1240520751, `RNS_PRIME_BITS'd1890021710, `RNS_PRIME_BITS'd1714689635, `RNS_PRIME_BITS'd1837319933, `RNS_PRIME_BITS'd147430926},
			'{`RNS_PRIME_BITS'd71, `RNS_PRIME_BITS'd1565957828, `RNS_PRIME_BITS'd1991286256, `RNS_PRIME_BITS'd1270441730, `RNS_PRIME_BITS'd219503422, `RNS_PRIME_BITS'd1691331767, `RNS_PRIME_BITS'd688839512, `RNS_PRIME_BITS'd1229997577, `RNS_PRIME_BITS'd892592915, `RNS_PRIME_BITS'd1126581775, `RNS_PRIME_BITS'd585949741},
			'{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd1369063276, `RNS_PRIME_BITS'd866358980, `RNS_PRIME_BITS'd549408617, `RNS_PRIME_BITS'd1586899871, `RNS_PRIME_BITS'd1764138862, `RNS_PRIME_BITS'd1769630713, `RNS_PRIME_BITS'd851065441, `RNS_PRIME_BITS'd1662313367, `RNS_PRIME_BITS'd439504921, `RNS_PRIME_BITS'd282411524},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1814409216, `RNS_PRIME_BITS'd2057101126, `RNS_PRIME_BITS'd2128492248, `RNS_PRIME_BITS'd303838695, `RNS_PRIME_BITS'd129755776, `RNS_PRIME_BITS'd1017090795, `RNS_PRIME_BITS'd1309600589, `RNS_PRIME_BITS'd2097196418, `RNS_PRIME_BITS'd821960401, `RNS_PRIME_BITS'd264648777},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd1291810513, `RNS_PRIME_BITS'd1788845809, `RNS_PRIME_BITS'd965489018, `RNS_PRIME_BITS'd1997490397, `RNS_PRIME_BITS'd1757305924, `RNS_PRIME_BITS'd730207898, `RNS_PRIME_BITS'd456676942, `RNS_PRIME_BITS'd925828563, `RNS_PRIME_BITS'd2145376410, `RNS_PRIME_BITS'd1191714465},
			'{`RNS_PRIME_BITS'd180, `RNS_PRIME_BITS'd735141042, `RNS_PRIME_BITS'd851750904, `RNS_PRIME_BITS'd1085835858, `RNS_PRIME_BITS'd924131462, `RNS_PRIME_BITS'd306122047, `RNS_PRIME_BITS'd952484028, `RNS_PRIME_BITS'd708601895, `RNS_PRIME_BITS'd216086993, `RNS_PRIME_BITS'd940275477, `RNS_PRIME_BITS'd985099135},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd1267726868, `RNS_PRIME_BITS'd212466890, `RNS_PRIME_BITS'd68827466, `RNS_PRIME_BITS'd432568065, `RNS_PRIME_BITS'd949705862, `RNS_PRIME_BITS'd614829181, `RNS_PRIME_BITS'd341331633, `RNS_PRIME_BITS'd1340500112, `RNS_PRIME_BITS'd1354222277, `RNS_PRIME_BITS'd2086545886},
			'{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd412012672, `RNS_PRIME_BITS'd403005071, `RNS_PRIME_BITS'd972335272, `RNS_PRIME_BITS'd484522196, `RNS_PRIME_BITS'd1645429793, `RNS_PRIME_BITS'd2044104438, `RNS_PRIME_BITS'd881615171, `RNS_PRIME_BITS'd1234306395, `RNS_PRIME_BITS'd884639471, `RNS_PRIME_BITS'd1204387166},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1187311937, `RNS_PRIME_BITS'd1797626571, `RNS_PRIME_BITS'd629943944, `RNS_PRIME_BITS'd663712091, `RNS_PRIME_BITS'd1139796089, `RNS_PRIME_BITS'd1801739604, `RNS_PRIME_BITS'd1760801499, `RNS_PRIME_BITS'd926130983, `RNS_PRIME_BITS'd334902519, `RNS_PRIME_BITS'd974871474},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd1403003378, `RNS_PRIME_BITS'd724869192, `RNS_PRIME_BITS'd1389720451, `RNS_PRIME_BITS'd791535971, `RNS_PRIME_BITS'd1804555789, `RNS_PRIME_BITS'd1345067108, `RNS_PRIME_BITS'd1359888201, `RNS_PRIME_BITS'd579464848, `RNS_PRIME_BITS'd530521964, `RNS_PRIME_BITS'd1682479150},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1650551055, `RNS_PRIME_BITS'd887901777, `RNS_PRIME_BITS'd1945950614, `RNS_PRIME_BITS'd2038485919, `RNS_PRIME_BITS'd284978867, `RNS_PRIME_BITS'd809347126, `RNS_PRIME_BITS'd1567239060, `RNS_PRIME_BITS'd1383197789, `RNS_PRIME_BITS'd2045854944, `RNS_PRIME_BITS'd1962765131},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1246832992, `RNS_PRIME_BITS'd1190200593, `RNS_PRIME_BITS'd273918758, `RNS_PRIME_BITS'd756362185, `RNS_PRIME_BITS'd1150296081, `RNS_PRIME_BITS'd1659384456, `RNS_PRIME_BITS'd1418731572, `RNS_PRIME_BITS'd584870409, `RNS_PRIME_BITS'd701478225, `RNS_PRIME_BITS'd383675401},
			'{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd1003181354, `RNS_PRIME_BITS'd157945717, `RNS_PRIME_BITS'd156595136, `RNS_PRIME_BITS'd150346886, `RNS_PRIME_BITS'd1871450636, `RNS_PRIME_BITS'd1406210475, `RNS_PRIME_BITS'd1630073408, `RNS_PRIME_BITS'd366352988, `RNS_PRIME_BITS'd378370534, `RNS_PRIME_BITS'd1722625291},
			'{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd965365729, `RNS_PRIME_BITS'd1162800917, `RNS_PRIME_BITS'd1149462843, `RNS_PRIME_BITS'd497816576, `RNS_PRIME_BITS'd1314336627, `RNS_PRIME_BITS'd482506731, `RNS_PRIME_BITS'd1965700036, `RNS_PRIME_BITS'd1804534115, `RNS_PRIME_BITS'd802263164, `RNS_PRIME_BITS'd392567835},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd61794611, `RNS_PRIME_BITS'd1595983014, `RNS_PRIME_BITS'd231721729, `RNS_PRIME_BITS'd1951902849, `RNS_PRIME_BITS'd1491035072, `RNS_PRIME_BITS'd379428464, `RNS_PRIME_BITS'd773445703, `RNS_PRIME_BITS'd1097754701, `RNS_PRIME_BITS'd552942801, `RNS_PRIME_BITS'd197727513},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd134307229, `RNS_PRIME_BITS'd1179606513, `RNS_PRIME_BITS'd337060499, `RNS_PRIME_BITS'd1118904309, `RNS_PRIME_BITS'd777115150, `RNS_PRIME_BITS'd686053284, `RNS_PRIME_BITS'd1159971279, `RNS_PRIME_BITS'd278627732, `RNS_PRIME_BITS'd245787442, `RNS_PRIME_BITS'd210286371},
			'{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd2097541729, `RNS_PRIME_BITS'd837196778, `RNS_PRIME_BITS'd43312718, `RNS_PRIME_BITS'd1683479087, `RNS_PRIME_BITS'd1488004477, `RNS_PRIME_BITS'd837717797, `RNS_PRIME_BITS'd1353154391, `RNS_PRIME_BITS'd523716189, `RNS_PRIME_BITS'd183205047, `RNS_PRIME_BITS'd918175577},
			'{`RNS_PRIME_BITS'd230, `RNS_PRIME_BITS'd1729028447, `RNS_PRIME_BITS'd500733241, `RNS_PRIME_BITS'd497230928, `RNS_PRIME_BITS'd2042759947, `RNS_PRIME_BITS'd1486225929, `RNS_PRIME_BITS'd328030269, `RNS_PRIME_BITS'd575940372, `RNS_PRIME_BITS'd1572789866, `RNS_PRIME_BITS'd2006900132, `RNS_PRIME_BITS'd959540451},
			'{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd783621845, `RNS_PRIME_BITS'd923212497, `RNS_PRIME_BITS'd1649151263, `RNS_PRIME_BITS'd1462535597, `RNS_PRIME_BITS'd20338309, `RNS_PRIME_BITS'd716657530, `RNS_PRIME_BITS'd1198576395, `RNS_PRIME_BITS'd2045697702, `RNS_PRIME_BITS'd73149826, `RNS_PRIME_BITS'd550536932},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd863875597, `RNS_PRIME_BITS'd234952816, `RNS_PRIME_BITS'd2039384472, `RNS_PRIME_BITS'd213212807, `RNS_PRIME_BITS'd1671205382, `RNS_PRIME_BITS'd2024740297, `RNS_PRIME_BITS'd43785035, `RNS_PRIME_BITS'd275788902, `RNS_PRIME_BITS'd2050658408, `RNS_PRIME_BITS'd389587171}
		},
		'{
			'{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd1067967450, `RNS_PRIME_BITS'd675732697, `RNS_PRIME_BITS'd285260077, `RNS_PRIME_BITS'd211597274, `RNS_PRIME_BITS'd356179392, `RNS_PRIME_BITS'd5168544, `RNS_PRIME_BITS'd172599261, `RNS_PRIME_BITS'd1981595514, `RNS_PRIME_BITS'd896632515, `RNS_PRIME_BITS'd882599369},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd494571271, `RNS_PRIME_BITS'd848912063, `RNS_PRIME_BITS'd281093768, `RNS_PRIME_BITS'd1164137236, `RNS_PRIME_BITS'd888581727, `RNS_PRIME_BITS'd401713180, `RNS_PRIME_BITS'd1849215982, `RNS_PRIME_BITS'd2100403981, `RNS_PRIME_BITS'd1364422947, `RNS_PRIME_BITS'd883132465},
			'{`RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd1403334048, `RNS_PRIME_BITS'd1614446436, `RNS_PRIME_BITS'd1715723218, `RNS_PRIME_BITS'd186003800, `RNS_PRIME_BITS'd745377445, `RNS_PRIME_BITS'd2116159705, `RNS_PRIME_BITS'd228704680, `RNS_PRIME_BITS'd941252873, `RNS_PRIME_BITS'd289757708, `RNS_PRIME_BITS'd2056107614},
			'{`RNS_PRIME_BITS'd238, `RNS_PRIME_BITS'd2089783162, `RNS_PRIME_BITS'd931998078, `RNS_PRIME_BITS'd904804499, `RNS_PRIME_BITS'd681754481, `RNS_PRIME_BITS'd996063947, `RNS_PRIME_BITS'd238678435, `RNS_PRIME_BITS'd648826075, `RNS_PRIME_BITS'd2021260666, `RNS_PRIME_BITS'd1744141181, `RNS_PRIME_BITS'd313216727},
			'{`RNS_PRIME_BITS'd69, `RNS_PRIME_BITS'd539923165, `RNS_PRIME_BITS'd1359636762, `RNS_PRIME_BITS'd1416690289, `RNS_PRIME_BITS'd313170236, `RNS_PRIME_BITS'd118353331, `RNS_PRIME_BITS'd1172645383, `RNS_PRIME_BITS'd187814541, `RNS_PRIME_BITS'd1469571860, `RNS_PRIME_BITS'd1683736740, `RNS_PRIME_BITS'd591023516},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd698607113, `RNS_PRIME_BITS'd1923156466, `RNS_PRIME_BITS'd93704250, `RNS_PRIME_BITS'd1998040195, `RNS_PRIME_BITS'd301103714, `RNS_PRIME_BITS'd1540642046, `RNS_PRIME_BITS'd2028042048, `RNS_PRIME_BITS'd235170380, `RNS_PRIME_BITS'd1408907703, `RNS_PRIME_BITS'd246115850},
			'{`RNS_PRIME_BITS'd254, `RNS_PRIME_BITS'd247114824, `RNS_PRIME_BITS'd1885756864, `RNS_PRIME_BITS'd1355258057, `RNS_PRIME_BITS'd2025355597, `RNS_PRIME_BITS'd1662237327, `RNS_PRIME_BITS'd1918337825, `RNS_PRIME_BITS'd2018546115, `RNS_PRIME_BITS'd92369285, `RNS_PRIME_BITS'd1799365468, `RNS_PRIME_BITS'd644177493},
			'{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd168148498, `RNS_PRIME_BITS'd1779721865, `RNS_PRIME_BITS'd163033101, `RNS_PRIME_BITS'd1750869053, `RNS_PRIME_BITS'd412490649, `RNS_PRIME_BITS'd1067412783, `RNS_PRIME_BITS'd882893238, `RNS_PRIME_BITS'd913254015, `RNS_PRIME_BITS'd426827509, `RNS_PRIME_BITS'd1838666343},
			'{`RNS_PRIME_BITS'd86, `RNS_PRIME_BITS'd1418655377, `RNS_PRIME_BITS'd1434842563, `RNS_PRIME_BITS'd906829818, `RNS_PRIME_BITS'd65315593, `RNS_PRIME_BITS'd1611013607, `RNS_PRIME_BITS'd1299149177, `RNS_PRIME_BITS'd1548711771, `RNS_PRIME_BITS'd1816244228, `RNS_PRIME_BITS'd236216235, `RNS_PRIME_BITS'd584872486},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1321485482, `RNS_PRIME_BITS'd496530283, `RNS_PRIME_BITS'd86675899, `RNS_PRIME_BITS'd2009889669, `RNS_PRIME_BITS'd1113546686, `RNS_PRIME_BITS'd1395096989, `RNS_PRIME_BITS'd319000608, `RNS_PRIME_BITS'd584859445, `RNS_PRIME_BITS'd1664373406, `RNS_PRIME_BITS'd462340276},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd313432471, `RNS_PRIME_BITS'd1652774172, `RNS_PRIME_BITS'd1730563623, `RNS_PRIME_BITS'd961415862, `RNS_PRIME_BITS'd1798629476, `RNS_PRIME_BITS'd1334988223, `RNS_PRIME_BITS'd623321868, `RNS_PRIME_BITS'd742552904, `RNS_PRIME_BITS'd327409473, `RNS_PRIME_BITS'd10524014},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1997226064, `RNS_PRIME_BITS'd2126888162, `RNS_PRIME_BITS'd1497131613, `RNS_PRIME_BITS'd186429585, `RNS_PRIME_BITS'd1343011348, `RNS_PRIME_BITS'd691218174, `RNS_PRIME_BITS'd964010165, `RNS_PRIME_BITS'd1428422582, `RNS_PRIME_BITS'd553229454, `RNS_PRIME_BITS'd256834528},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd1127700632, `RNS_PRIME_BITS'd563750069, `RNS_PRIME_BITS'd1871691342, `RNS_PRIME_BITS'd1831336670, `RNS_PRIME_BITS'd1153224354, `RNS_PRIME_BITS'd1504472071, `RNS_PRIME_BITS'd947145196, `RNS_PRIME_BITS'd82206977, `RNS_PRIME_BITS'd730151309, `RNS_PRIME_BITS'd2015009057},
			'{`RNS_PRIME_BITS'd165, `RNS_PRIME_BITS'd1299503992, `RNS_PRIME_BITS'd6606655, `RNS_PRIME_BITS'd157760184, `RNS_PRIME_BITS'd1456084820, `RNS_PRIME_BITS'd635875504, `RNS_PRIME_BITS'd1538081271, `RNS_PRIME_BITS'd1175658035, `RNS_PRIME_BITS'd762338298, `RNS_PRIME_BITS'd58928530, `RNS_PRIME_BITS'd333743840},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1207226092, `RNS_PRIME_BITS'd1764976255, `RNS_PRIME_BITS'd459774286, `RNS_PRIME_BITS'd845164119, `RNS_PRIME_BITS'd1569932331, `RNS_PRIME_BITS'd1441713672, `RNS_PRIME_BITS'd2073776679, `RNS_PRIME_BITS'd1490777854, `RNS_PRIME_BITS'd1480687151, `RNS_PRIME_BITS'd480160357},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd1415338265, `RNS_PRIME_BITS'd1535184560, `RNS_PRIME_BITS'd68265057, `RNS_PRIME_BITS'd2029515296, `RNS_PRIME_BITS'd2022470597, `RNS_PRIME_BITS'd1238192738, `RNS_PRIME_BITS'd1914388633, `RNS_PRIME_BITS'd335004962, `RNS_PRIME_BITS'd1519309713, `RNS_PRIME_BITS'd791907525},
			'{`RNS_PRIME_BITS'd180, `RNS_PRIME_BITS'd270466085, `RNS_PRIME_BITS'd1813499936, `RNS_PRIME_BITS'd516496983, `RNS_PRIME_BITS'd805615709, `RNS_PRIME_BITS'd1502313803, `RNS_PRIME_BITS'd1437411443, `RNS_PRIME_BITS'd1470714454, `RNS_PRIME_BITS'd1251502395, `RNS_PRIME_BITS'd716676739, `RNS_PRIME_BITS'd1407775533},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd1400909828, `RNS_PRIME_BITS'd1593088348, `RNS_PRIME_BITS'd264973178, `RNS_PRIME_BITS'd1320671372, `RNS_PRIME_BITS'd7727565, `RNS_PRIME_BITS'd16488147, `RNS_PRIME_BITS'd267778832, `RNS_PRIME_BITS'd378964322, `RNS_PRIME_BITS'd1937646163, `RNS_PRIME_BITS'd677018325},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd1060673046, `RNS_PRIME_BITS'd93760284, `RNS_PRIME_BITS'd881571602, `RNS_PRIME_BITS'd1129869602, `RNS_PRIME_BITS'd285420527, `RNS_PRIME_BITS'd2049375072, `RNS_PRIME_BITS'd1486306390, `RNS_PRIME_BITS'd1113906822, `RNS_PRIME_BITS'd1673993456, `RNS_PRIME_BITS'd413684776},
			'{`RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd225567157, `RNS_PRIME_BITS'd1150933316, `RNS_PRIME_BITS'd1348726102, `RNS_PRIME_BITS'd951477055, `RNS_PRIME_BITS'd1285405322, `RNS_PRIME_BITS'd960951667, `RNS_PRIME_BITS'd1071532018, `RNS_PRIME_BITS'd335586659, `RNS_PRIME_BITS'd97839328, `RNS_PRIME_BITS'd1829876398},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1667069791, `RNS_PRIME_BITS'd143301128, `RNS_PRIME_BITS'd400947515, `RNS_PRIME_BITS'd1652187910, `RNS_PRIME_BITS'd1260359150, `RNS_PRIME_BITS'd1967064846, `RNS_PRIME_BITS'd1688430528, `RNS_PRIME_BITS'd382625687, `RNS_PRIME_BITS'd1249467709, `RNS_PRIME_BITS'd1324008597},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd2110313560, `RNS_PRIME_BITS'd266828444, `RNS_PRIME_BITS'd930691400, `RNS_PRIME_BITS'd49431275, `RNS_PRIME_BITS'd70063156, `RNS_PRIME_BITS'd1990232920, `RNS_PRIME_BITS'd42523414, `RNS_PRIME_BITS'd552243080, `RNS_PRIME_BITS'd366803284, `RNS_PRIME_BITS'd429064310},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd2070519602, `RNS_PRIME_BITS'd2006336897, `RNS_PRIME_BITS'd1425947176, `RNS_PRIME_BITS'd539316340, `RNS_PRIME_BITS'd899544233, `RNS_PRIME_BITS'd658118695, `RNS_PRIME_BITS'd607144528, `RNS_PRIME_BITS'd2008700509, `RNS_PRIME_BITS'd734229588, `RNS_PRIME_BITS'd2006166632},
			'{`RNS_PRIME_BITS'd151, `RNS_PRIME_BITS'd918783669, `RNS_PRIME_BITS'd1716406138, `RNS_PRIME_BITS'd1264401040, `RNS_PRIME_BITS'd1969206537, `RNS_PRIME_BITS'd1943134679, `RNS_PRIME_BITS'd942805112, `RNS_PRIME_BITS'd535657216, `RNS_PRIME_BITS'd2094576006, `RNS_PRIME_BITS'd1461039985, `RNS_PRIME_BITS'd870620432},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd1275200574, `RNS_PRIME_BITS'd1576469921, `RNS_PRIME_BITS'd605897511, `RNS_PRIME_BITS'd754190940, `RNS_PRIME_BITS'd1509128080, `RNS_PRIME_BITS'd268145989, `RNS_PRIME_BITS'd63011650, `RNS_PRIME_BITS'd306276452, `RNS_PRIME_BITS'd1514111611, `RNS_PRIME_BITS'd68021235},
			'{`RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd604048473, `RNS_PRIME_BITS'd274346655, `RNS_PRIME_BITS'd935627088, `RNS_PRIME_BITS'd249792907, `RNS_PRIME_BITS'd650195281, `RNS_PRIME_BITS'd495165067, `RNS_PRIME_BITS'd2067534261, `RNS_PRIME_BITS'd368912264, `RNS_PRIME_BITS'd878468279, `RNS_PRIME_BITS'd933620386},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd691638126, `RNS_PRIME_BITS'd1197322048, `RNS_PRIME_BITS'd300875213, `RNS_PRIME_BITS'd726320777, `RNS_PRIME_BITS'd2130796484, `RNS_PRIME_BITS'd2055170488, `RNS_PRIME_BITS'd1066034117, `RNS_PRIME_BITS'd1838737075, `RNS_PRIME_BITS'd431217898, `RNS_PRIME_BITS'd1610523404},
			'{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd118022012, `RNS_PRIME_BITS'd1901054774, `RNS_PRIME_BITS'd1599345044, `RNS_PRIME_BITS'd1409990469, `RNS_PRIME_BITS'd1457658226, `RNS_PRIME_BITS'd99118029, `RNS_PRIME_BITS'd1838876321, `RNS_PRIME_BITS'd1950000656, `RNS_PRIME_BITS'd1196799089, `RNS_PRIME_BITS'd1835051861},
			'{`RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd277322771, `RNS_PRIME_BITS'd2139913820, `RNS_PRIME_BITS'd386239283, `RNS_PRIME_BITS'd310451681, `RNS_PRIME_BITS'd537621489, `RNS_PRIME_BITS'd1653506491, `RNS_PRIME_BITS'd66332358, `RNS_PRIME_BITS'd1429079204, `RNS_PRIME_BITS'd1993987391, `RNS_PRIME_BITS'd1586304399},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1060247167, `RNS_PRIME_BITS'd988419822, `RNS_PRIME_BITS'd260225606, `RNS_PRIME_BITS'd419858562, `RNS_PRIME_BITS'd1892324948, `RNS_PRIME_BITS'd988930034, `RNS_PRIME_BITS'd1128150710, `RNS_PRIME_BITS'd1228427638, `RNS_PRIME_BITS'd1429234976, `RNS_PRIME_BITS'd1334273445},
			'{`RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd160906088, `RNS_PRIME_BITS'd1962814803, `RNS_PRIME_BITS'd985261670, `RNS_PRIME_BITS'd489611319, `RNS_PRIME_BITS'd1931406893, `RNS_PRIME_BITS'd11535858, `RNS_PRIME_BITS'd352461250, `RNS_PRIME_BITS'd111419101, `RNS_PRIME_BITS'd1085692448, `RNS_PRIME_BITS'd1508855799},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd1644120659, `RNS_PRIME_BITS'd1639487671, `RNS_PRIME_BITS'd187543081, `RNS_PRIME_BITS'd1407020219, `RNS_PRIME_BITS'd2042099914, `RNS_PRIME_BITS'd1640200972, `RNS_PRIME_BITS'd1592373564, `RNS_PRIME_BITS'd2075249453, `RNS_PRIME_BITS'd1398795032, `RNS_PRIME_BITS'd492311315},
			'{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd122080978, `RNS_PRIME_BITS'd349231878, `RNS_PRIME_BITS'd1720609214, `RNS_PRIME_BITS'd296981313, `RNS_PRIME_BITS'd928252864, `RNS_PRIME_BITS'd275594869, `RNS_PRIME_BITS'd907984584, `RNS_PRIME_BITS'd1780331253, `RNS_PRIME_BITS'd2132043053, `RNS_PRIME_BITS'd572035538},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd2127353293, `RNS_PRIME_BITS'd1874836084, `RNS_PRIME_BITS'd1841950617, `RNS_PRIME_BITS'd1219006834, `RNS_PRIME_BITS'd1931855365, `RNS_PRIME_BITS'd618657970, `RNS_PRIME_BITS'd763750858, `RNS_PRIME_BITS'd84214321, `RNS_PRIME_BITS'd1640291024, `RNS_PRIME_BITS'd2135149865},
			'{`RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd2115374764, `RNS_PRIME_BITS'd818025809, `RNS_PRIME_BITS'd1934459606, `RNS_PRIME_BITS'd447984242, `RNS_PRIME_BITS'd235341351, `RNS_PRIME_BITS'd1070703554, `RNS_PRIME_BITS'd951168761, `RNS_PRIME_BITS'd8847818, `RNS_PRIME_BITS'd790348726, `RNS_PRIME_BITS'd72248052},
			'{`RNS_PRIME_BITS'd14, `RNS_PRIME_BITS'd51203610, `RNS_PRIME_BITS'd779312764, `RNS_PRIME_BITS'd181464161, `RNS_PRIME_BITS'd1255260337, `RNS_PRIME_BITS'd1097830735, `RNS_PRIME_BITS'd803072662, `RNS_PRIME_BITS'd1245631061, `RNS_PRIME_BITS'd1419670714, `RNS_PRIME_BITS'd2113079321, `RNS_PRIME_BITS'd891214438},
			'{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd295210506, `RNS_PRIME_BITS'd613460651, `RNS_PRIME_BITS'd1629762888, `RNS_PRIME_BITS'd1013888645, `RNS_PRIME_BITS'd1799534366, `RNS_PRIME_BITS'd1251033017, `RNS_PRIME_BITS'd115531826, `RNS_PRIME_BITS'd1883753837, `RNS_PRIME_BITS'd757756391, `RNS_PRIME_BITS'd800908932},
			'{`RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd617168222, `RNS_PRIME_BITS'd209693244, `RNS_PRIME_BITS'd76586956, `RNS_PRIME_BITS'd817491829, `RNS_PRIME_BITS'd1439585057, `RNS_PRIME_BITS'd747735522, `RNS_PRIME_BITS'd1873129710, `RNS_PRIME_BITS'd1949723305, `RNS_PRIME_BITS'd1275286453, `RNS_PRIME_BITS'd651620233},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1953617632, `RNS_PRIME_BITS'd197587191, `RNS_PRIME_BITS'd1338244205, `RNS_PRIME_BITS'd2014869717, `RNS_PRIME_BITS'd1320483227, `RNS_PRIME_BITS'd375250902, `RNS_PRIME_BITS'd835035460, `RNS_PRIME_BITS'd1228044869, `RNS_PRIME_BITS'd1221908686, `RNS_PRIME_BITS'd1203053042},
			'{`RNS_PRIME_BITS'd172, `RNS_PRIME_BITS'd1041254052, `RNS_PRIME_BITS'd986463267, `RNS_PRIME_BITS'd10583415, `RNS_PRIME_BITS'd119878454, `RNS_PRIME_BITS'd1185264846, `RNS_PRIME_BITS'd1685734034, `RNS_PRIME_BITS'd1485198765, `RNS_PRIME_BITS'd376085577, `RNS_PRIME_BITS'd1412499985, `RNS_PRIME_BITS'd897885584},
			'{`RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd1611160931, `RNS_PRIME_BITS'd315106836, `RNS_PRIME_BITS'd1078281798, `RNS_PRIME_BITS'd1475020536, `RNS_PRIME_BITS'd971556876, `RNS_PRIME_BITS'd1917257848, `RNS_PRIME_BITS'd1367011360, `RNS_PRIME_BITS'd1050002796, `RNS_PRIME_BITS'd1471875740, `RNS_PRIME_BITS'd4991108},
			'{`RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd591833009, `RNS_PRIME_BITS'd2142546002, `RNS_PRIME_BITS'd294953032, `RNS_PRIME_BITS'd1168947880, `RNS_PRIME_BITS'd253649657, `RNS_PRIME_BITS'd1443161497, `RNS_PRIME_BITS'd967454043, `RNS_PRIME_BITS'd1267149936, `RNS_PRIME_BITS'd1502308518, `RNS_PRIME_BITS'd1895894885},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd780940226, `RNS_PRIME_BITS'd1379790540, `RNS_PRIME_BITS'd1855570864, `RNS_PRIME_BITS'd2123487539, `RNS_PRIME_BITS'd1062527381, `RNS_PRIME_BITS'd1376565020, `RNS_PRIME_BITS'd915807088, `RNS_PRIME_BITS'd1115970748, `RNS_PRIME_BITS'd1073957144, `RNS_PRIME_BITS'd1958202362},
			'{`RNS_PRIME_BITS'd40, `RNS_PRIME_BITS'd1267188117, `RNS_PRIME_BITS'd2145349923, `RNS_PRIME_BITS'd1936490391, `RNS_PRIME_BITS'd1058856382, `RNS_PRIME_BITS'd610173993, `RNS_PRIME_BITS'd1652300176, `RNS_PRIME_BITS'd1280495219, `RNS_PRIME_BITS'd318210620, `RNS_PRIME_BITS'd632551175, `RNS_PRIME_BITS'd1624172372},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd2057715565, `RNS_PRIME_BITS'd904840892, `RNS_PRIME_BITS'd516504888, `RNS_PRIME_BITS'd95757193, `RNS_PRIME_BITS'd526953189, `RNS_PRIME_BITS'd2105672120, `RNS_PRIME_BITS'd1109966926, `RNS_PRIME_BITS'd1723621631, `RNS_PRIME_BITS'd630649480, `RNS_PRIME_BITS'd1335250529},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd240819087, `RNS_PRIME_BITS'd2067319700, `RNS_PRIME_BITS'd849702492, `RNS_PRIME_BITS'd1267832862, `RNS_PRIME_BITS'd1006088918, `RNS_PRIME_BITS'd78579015, `RNS_PRIME_BITS'd70207309, `RNS_PRIME_BITS'd1041481304, `RNS_PRIME_BITS'd1515555665, `RNS_PRIME_BITS'd820639890},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd147998877, `RNS_PRIME_BITS'd2059406843, `RNS_PRIME_BITS'd1565814915, `RNS_PRIME_BITS'd1194590728, `RNS_PRIME_BITS'd1551704052, `RNS_PRIME_BITS'd1725600033, `RNS_PRIME_BITS'd1690430718, `RNS_PRIME_BITS'd2041902494, `RNS_PRIME_BITS'd1673675130, `RNS_PRIME_BITS'd697118648},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1095379058, `RNS_PRIME_BITS'd21572574, `RNS_PRIME_BITS'd331261161, `RNS_PRIME_BITS'd191113905, `RNS_PRIME_BITS'd2138028339, `RNS_PRIME_BITS'd483581508, `RNS_PRIME_BITS'd499221240, `RNS_PRIME_BITS'd1418508038, `RNS_PRIME_BITS'd2076061237, `RNS_PRIME_BITS'd209377478},
			'{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd749385872, `RNS_PRIME_BITS'd905380176, `RNS_PRIME_BITS'd1425541696, `RNS_PRIME_BITS'd483749878, `RNS_PRIME_BITS'd896078943, `RNS_PRIME_BITS'd894009874, `RNS_PRIME_BITS'd1815459850, `RNS_PRIME_BITS'd1404354122, `RNS_PRIME_BITS'd1075537443, `RNS_PRIME_BITS'd1025765602},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd233632476, `RNS_PRIME_BITS'd1989913779, `RNS_PRIME_BITS'd2100066691, `RNS_PRIME_BITS'd759252062, `RNS_PRIME_BITS'd1650554059, `RNS_PRIME_BITS'd2110391080, `RNS_PRIME_BITS'd67355135, `RNS_PRIME_BITS'd1866504371, `RNS_PRIME_BITS'd1852695689, `RNS_PRIME_BITS'd1018395345},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd922841961, `RNS_PRIME_BITS'd1511303724, `RNS_PRIME_BITS'd1289329097, `RNS_PRIME_BITS'd1119462188, `RNS_PRIME_BITS'd2038222520, `RNS_PRIME_BITS'd991018652, `RNS_PRIME_BITS'd697505123, `RNS_PRIME_BITS'd659004716, `RNS_PRIME_BITS'd364533845, `RNS_PRIME_BITS'd304350246},
			'{`RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd859696064, `RNS_PRIME_BITS'd456771337, `RNS_PRIME_BITS'd656267601, `RNS_PRIME_BITS'd2113085009, `RNS_PRIME_BITS'd518265863, `RNS_PRIME_BITS'd1927260746, `RNS_PRIME_BITS'd388858847, `RNS_PRIME_BITS'd2019814068, `RNS_PRIME_BITS'd43229109, `RNS_PRIME_BITS'd1777857592},
			'{`RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd1878229338, `RNS_PRIME_BITS'd1369986087, `RNS_PRIME_BITS'd1608717247, `RNS_PRIME_BITS'd1109489895, `RNS_PRIME_BITS'd545538833, `RNS_PRIME_BITS'd26931056, `RNS_PRIME_BITS'd60665634, `RNS_PRIME_BITS'd986527215, `RNS_PRIME_BITS'd134715290, `RNS_PRIME_BITS'd492164241},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1938167985, `RNS_PRIME_BITS'd654402852, `RNS_PRIME_BITS'd321126528, `RNS_PRIME_BITS'd675752526, `RNS_PRIME_BITS'd75690734, `RNS_PRIME_BITS'd1149458368, `RNS_PRIME_BITS'd932761650, `RNS_PRIME_BITS'd793531701, `RNS_PRIME_BITS'd641447625, `RNS_PRIME_BITS'd1199478854},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd602626029, `RNS_PRIME_BITS'd223175660, `RNS_PRIME_BITS'd291480216, `RNS_PRIME_BITS'd1352476065, `RNS_PRIME_BITS'd1130812134, `RNS_PRIME_BITS'd802021040, `RNS_PRIME_BITS'd1361582433, `RNS_PRIME_BITS'd1811086133, `RNS_PRIME_BITS'd1320228919, `RNS_PRIME_BITS'd1058731684},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1308571167, `RNS_PRIME_BITS'd625567877, `RNS_PRIME_BITS'd1766051342, `RNS_PRIME_BITS'd715705132, `RNS_PRIME_BITS'd1091433812, `RNS_PRIME_BITS'd504319132, `RNS_PRIME_BITS'd1707298107, `RNS_PRIME_BITS'd914841515, `RNS_PRIME_BITS'd324605966, `RNS_PRIME_BITS'd1196904792},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd1112722181, `RNS_PRIME_BITS'd1605334825, `RNS_PRIME_BITS'd2068975932, `RNS_PRIME_BITS'd254648932, `RNS_PRIME_BITS'd221006334, `RNS_PRIME_BITS'd1984617920, `RNS_PRIME_BITS'd114130997, `RNS_PRIME_BITS'd2039511045, `RNS_PRIME_BITS'd616730191, `RNS_PRIME_BITS'd1056137745},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd369541506, `RNS_PRIME_BITS'd756949738, `RNS_PRIME_BITS'd1356851945, `RNS_PRIME_BITS'd577910903, `RNS_PRIME_BITS'd1680265387, `RNS_PRIME_BITS'd992944381, `RNS_PRIME_BITS'd218235379, `RNS_PRIME_BITS'd1933797353, `RNS_PRIME_BITS'd628968090, `RNS_PRIME_BITS'd407040416},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd1748446179, `RNS_PRIME_BITS'd612973495, `RNS_PRIME_BITS'd1201231948, `RNS_PRIME_BITS'd1509257284, `RNS_PRIME_BITS'd1084166834, `RNS_PRIME_BITS'd1488191624, `RNS_PRIME_BITS'd1115592509, `RNS_PRIME_BITS'd81680366, `RNS_PRIME_BITS'd862173632, `RNS_PRIME_BITS'd1236733456},
			'{`RNS_PRIME_BITS'd110, `RNS_PRIME_BITS'd1727847452, `RNS_PRIME_BITS'd672788045, `RNS_PRIME_BITS'd1073356003, `RNS_PRIME_BITS'd1096173568, `RNS_PRIME_BITS'd1287960388, `RNS_PRIME_BITS'd1258997834, `RNS_PRIME_BITS'd1559839525, `RNS_PRIME_BITS'd1989706008, `RNS_PRIME_BITS'd1175737772, `RNS_PRIME_BITS'd102948820},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd418280316, `RNS_PRIME_BITS'd1974754703, `RNS_PRIME_BITS'd601811378, `RNS_PRIME_BITS'd1987664443, `RNS_PRIME_BITS'd1116080339, `RNS_PRIME_BITS'd90847644, `RNS_PRIME_BITS'd1313983545, `RNS_PRIME_BITS'd853890271, `RNS_PRIME_BITS'd1683942945, `RNS_PRIME_BITS'd635828909},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd1253368156, `RNS_PRIME_BITS'd473373879, `RNS_PRIME_BITS'd1702552741, `RNS_PRIME_BITS'd1757484412, `RNS_PRIME_BITS'd1305867823, `RNS_PRIME_BITS'd1471919771, `RNS_PRIME_BITS'd1619545108, `RNS_PRIME_BITS'd310608863, `RNS_PRIME_BITS'd22257596, `RNS_PRIME_BITS'd3145909},
			'{`RNS_PRIME_BITS'd170, `RNS_PRIME_BITS'd1544681101, `RNS_PRIME_BITS'd1016777655, `RNS_PRIME_BITS'd1440875740, `RNS_PRIME_BITS'd776595645, `RNS_PRIME_BITS'd1356363439, `RNS_PRIME_BITS'd760592260, `RNS_PRIME_BITS'd1178031259, `RNS_PRIME_BITS'd245533048, `RNS_PRIME_BITS'd1905983377, `RNS_PRIME_BITS'd548821638},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd820919395, `RNS_PRIME_BITS'd275380717, `RNS_PRIME_BITS'd808900813, `RNS_PRIME_BITS'd1078522768, `RNS_PRIME_BITS'd418504500, `RNS_PRIME_BITS'd858808910, `RNS_PRIME_BITS'd1692385494, `RNS_PRIME_BITS'd1835367048, `RNS_PRIME_BITS'd1308743945, `RNS_PRIME_BITS'd1943976984}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd446123217, `RNS_PRIME_BITS'd1323396675, `RNS_PRIME_BITS'd1935258559, `RNS_PRIME_BITS'd1399662490, `RNS_PRIME_BITS'd329984314, `RNS_PRIME_BITS'd1464399932, `RNS_PRIME_BITS'd1847492473, `RNS_PRIME_BITS'd763010077, `RNS_PRIME_BITS'd336755007, `RNS_PRIME_BITS'd2074934023},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd181314914, `RNS_PRIME_BITS'd730550683, `RNS_PRIME_BITS'd590799953, `RNS_PRIME_BITS'd1391304750, `RNS_PRIME_BITS'd1784748612, `RNS_PRIME_BITS'd542418036, `RNS_PRIME_BITS'd1554795488, `RNS_PRIME_BITS'd476939289, `RNS_PRIME_BITS'd1344532666, `RNS_PRIME_BITS'd1837516088},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd1832094704, `RNS_PRIME_BITS'd898058095, `RNS_PRIME_BITS'd1657894406, `RNS_PRIME_BITS'd606652561, `RNS_PRIME_BITS'd652318589, `RNS_PRIME_BITS'd1894867456, `RNS_PRIME_BITS'd819942268, `RNS_PRIME_BITS'd1007924436, `RNS_PRIME_BITS'd100778698, `RNS_PRIME_BITS'd2114093760},
			'{`RNS_PRIME_BITS'd186, `RNS_PRIME_BITS'd1140453664, `RNS_PRIME_BITS'd552532672, `RNS_PRIME_BITS'd53854764, `RNS_PRIME_BITS'd1160048673, `RNS_PRIME_BITS'd1011258840, `RNS_PRIME_BITS'd2130818788, `RNS_PRIME_BITS'd959968451, `RNS_PRIME_BITS'd1010560246, `RNS_PRIME_BITS'd1579373700, `RNS_PRIME_BITS'd381113929},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd421776241, `RNS_PRIME_BITS'd1647165706, `RNS_PRIME_BITS'd226604321, `RNS_PRIME_BITS'd1101689684, `RNS_PRIME_BITS'd1655236857, `RNS_PRIME_BITS'd2052762805, `RNS_PRIME_BITS'd394591595, `RNS_PRIME_BITS'd1971440563, `RNS_PRIME_BITS'd1034278648, `RNS_PRIME_BITS'd192474969},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd241514381, `RNS_PRIME_BITS'd1839780618, `RNS_PRIME_BITS'd1906250892, `RNS_PRIME_BITS'd151896448, `RNS_PRIME_BITS'd631002911, `RNS_PRIME_BITS'd803892979, `RNS_PRIME_BITS'd1399314510, `RNS_PRIME_BITS'd578996934, `RNS_PRIME_BITS'd898718253, `RNS_PRIME_BITS'd1220080867},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd1402451192, `RNS_PRIME_BITS'd2143856328, `RNS_PRIME_BITS'd1048157940, `RNS_PRIME_BITS'd1215285180, `RNS_PRIME_BITS'd1182880489, `RNS_PRIME_BITS'd1059469751, `RNS_PRIME_BITS'd1416651122, `RNS_PRIME_BITS'd1809291300, `RNS_PRIME_BITS'd1683034035, `RNS_PRIME_BITS'd75639438},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd354677948, `RNS_PRIME_BITS'd1178262348, `RNS_PRIME_BITS'd274538589, `RNS_PRIME_BITS'd606236756, `RNS_PRIME_BITS'd946996215, `RNS_PRIME_BITS'd1429068824, `RNS_PRIME_BITS'd1766946659, `RNS_PRIME_BITS'd1614967309, `RNS_PRIME_BITS'd1291308780, `RNS_PRIME_BITS'd1503422289},
			'{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd1944796562, `RNS_PRIME_BITS'd1632194219, `RNS_PRIME_BITS'd951613702, `RNS_PRIME_BITS'd2136950431, `RNS_PRIME_BITS'd432935149, `RNS_PRIME_BITS'd838256977, `RNS_PRIME_BITS'd1097684140, `RNS_PRIME_BITS'd469517367, `RNS_PRIME_BITS'd48964568, `RNS_PRIME_BITS'd675150201},
			'{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd606360428, `RNS_PRIME_BITS'd26933662, `RNS_PRIME_BITS'd1247635058, `RNS_PRIME_BITS'd96587599, `RNS_PRIME_BITS'd801572975, `RNS_PRIME_BITS'd1603478709, `RNS_PRIME_BITS'd583982684, `RNS_PRIME_BITS'd50357986, `RNS_PRIME_BITS'd206003886, `RNS_PRIME_BITS'd1047061359},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd840502002, `RNS_PRIME_BITS'd113454960, `RNS_PRIME_BITS'd1621712631, `RNS_PRIME_BITS'd1974912430, `RNS_PRIME_BITS'd1543764931, `RNS_PRIME_BITS'd661901135, `RNS_PRIME_BITS'd80885482, `RNS_PRIME_BITS'd1702430063, `RNS_PRIME_BITS'd1431963600, `RNS_PRIME_BITS'd1622907753},
			'{`RNS_PRIME_BITS'd98, `RNS_PRIME_BITS'd809132347, `RNS_PRIME_BITS'd1228277704, `RNS_PRIME_BITS'd1183114276, `RNS_PRIME_BITS'd2026731153, `RNS_PRIME_BITS'd1871346371, `RNS_PRIME_BITS'd561135853, `RNS_PRIME_BITS'd1271266752, `RNS_PRIME_BITS'd322618879, `RNS_PRIME_BITS'd1799459013, `RNS_PRIME_BITS'd377527730},
			'{`RNS_PRIME_BITS'd148, `RNS_PRIME_BITS'd209778177, `RNS_PRIME_BITS'd102243267, `RNS_PRIME_BITS'd375170585, `RNS_PRIME_BITS'd1248178828, `RNS_PRIME_BITS'd828052166, `RNS_PRIME_BITS'd115772576, `RNS_PRIME_BITS'd404897407, `RNS_PRIME_BITS'd1559793278, `RNS_PRIME_BITS'd758791768, `RNS_PRIME_BITS'd1615235625},
			'{`RNS_PRIME_BITS'd220, `RNS_PRIME_BITS'd227153512, `RNS_PRIME_BITS'd998925361, `RNS_PRIME_BITS'd199323315, `RNS_PRIME_BITS'd1032937740, `RNS_PRIME_BITS'd713300169, `RNS_PRIME_BITS'd500667731, `RNS_PRIME_BITS'd2073212348, `RNS_PRIME_BITS'd644203539, `RNS_PRIME_BITS'd808287050, `RNS_PRIME_BITS'd1935753144},
			'{`RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd1946201092, `RNS_PRIME_BITS'd307476027, `RNS_PRIME_BITS'd2027606656, `RNS_PRIME_BITS'd997441507, `RNS_PRIME_BITS'd244210105, `RNS_PRIME_BITS'd1488660706, `RNS_PRIME_BITS'd1328063822, `RNS_PRIME_BITS'd611471256, `RNS_PRIME_BITS'd1667642719, `RNS_PRIME_BITS'd1524711549},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd51704212, `RNS_PRIME_BITS'd1565538672, `RNS_PRIME_BITS'd606356602, `RNS_PRIME_BITS'd1401724211, `RNS_PRIME_BITS'd63317993, `RNS_PRIME_BITS'd1262120564, `RNS_PRIME_BITS'd451431954, `RNS_PRIME_BITS'd1114647452, `RNS_PRIME_BITS'd1312683306, `RNS_PRIME_BITS'd628956923},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd1304736530, `RNS_PRIME_BITS'd2081634153, `RNS_PRIME_BITS'd1996645730, `RNS_PRIME_BITS'd1115369885, `RNS_PRIME_BITS'd1418938971, `RNS_PRIME_BITS'd257982187, `RNS_PRIME_BITS'd1600499315, `RNS_PRIME_BITS'd1203410259, `RNS_PRIME_BITS'd143322712, `RNS_PRIME_BITS'd1112918088},
			'{`RNS_PRIME_BITS'd32, `RNS_PRIME_BITS'd790255772, `RNS_PRIME_BITS'd1228429173, `RNS_PRIME_BITS'd1391630706, `RNS_PRIME_BITS'd684991964, `RNS_PRIME_BITS'd1653866924, `RNS_PRIME_BITS'd474757439, `RNS_PRIME_BITS'd6322318, `RNS_PRIME_BITS'd1084833115, `RNS_PRIME_BITS'd163201225, `RNS_PRIME_BITS'd496172726},
			'{`RNS_PRIME_BITS'd86, `RNS_PRIME_BITS'd1673758700, `RNS_PRIME_BITS'd477173065, `RNS_PRIME_BITS'd688799776, `RNS_PRIME_BITS'd1257328363, `RNS_PRIME_BITS'd240748995, `RNS_PRIME_BITS'd2136115906, `RNS_PRIME_BITS'd1539004075, `RNS_PRIME_BITS'd1465141720, `RNS_PRIME_BITS'd1772511746, `RNS_PRIME_BITS'd1549066184},
			'{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd44481972, `RNS_PRIME_BITS'd1555913310, `RNS_PRIME_BITS'd1075833146, `RNS_PRIME_BITS'd2000700666, `RNS_PRIME_BITS'd292540596, `RNS_PRIME_BITS'd350754168, `RNS_PRIME_BITS'd2065469460, `RNS_PRIME_BITS'd1669445538, `RNS_PRIME_BITS'd373261642, `RNS_PRIME_BITS'd559014197},
			'{`RNS_PRIME_BITS'd131, `RNS_PRIME_BITS'd966279963, `RNS_PRIME_BITS'd1366996084, `RNS_PRIME_BITS'd544943255, `RNS_PRIME_BITS'd932182029, `RNS_PRIME_BITS'd50723940, `RNS_PRIME_BITS'd430265713, `RNS_PRIME_BITS'd1784100541, `RNS_PRIME_BITS'd508608265, `RNS_PRIME_BITS'd774798266, `RNS_PRIME_BITS'd1779425731},
			'{`RNS_PRIME_BITS'd66, `RNS_PRIME_BITS'd934758331, `RNS_PRIME_BITS'd432095278, `RNS_PRIME_BITS'd65158339, `RNS_PRIME_BITS'd1795259491, `RNS_PRIME_BITS'd237252002, `RNS_PRIME_BITS'd419115706, `RNS_PRIME_BITS'd465487345, `RNS_PRIME_BITS'd746964093, `RNS_PRIME_BITS'd1536850680, `RNS_PRIME_BITS'd856724859},
			'{`RNS_PRIME_BITS'd15, `RNS_PRIME_BITS'd1788086089, `RNS_PRIME_BITS'd595354978, `RNS_PRIME_BITS'd247753740, `RNS_PRIME_BITS'd1327345325, `RNS_PRIME_BITS'd30187924, `RNS_PRIME_BITS'd1816609069, `RNS_PRIME_BITS'd457721345, `RNS_PRIME_BITS'd59312845, `RNS_PRIME_BITS'd625523152, `RNS_PRIME_BITS'd825215838},
			'{`RNS_PRIME_BITS'd230, `RNS_PRIME_BITS'd906817025, `RNS_PRIME_BITS'd909408754, `RNS_PRIME_BITS'd380619072, `RNS_PRIME_BITS'd668361610, `RNS_PRIME_BITS'd2017105975, `RNS_PRIME_BITS'd806162609, `RNS_PRIME_BITS'd19370997, `RNS_PRIME_BITS'd492255875, `RNS_PRIME_BITS'd181673825, `RNS_PRIME_BITS'd913329572},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd1289424245, `RNS_PRIME_BITS'd823755271, `RNS_PRIME_BITS'd1882375914, `RNS_PRIME_BITS'd2015267746, `RNS_PRIME_BITS'd898017303, `RNS_PRIME_BITS'd217971082, `RNS_PRIME_BITS'd443759553, `RNS_PRIME_BITS'd282748161, `RNS_PRIME_BITS'd1020553819, `RNS_PRIME_BITS'd747790430},
			'{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd1560406679, `RNS_PRIME_BITS'd323302168, `RNS_PRIME_BITS'd2051912762, `RNS_PRIME_BITS'd1992523004, `RNS_PRIME_BITS'd1620502651, `RNS_PRIME_BITS'd1920331572, `RNS_PRIME_BITS'd1816381894, `RNS_PRIME_BITS'd2104107064, `RNS_PRIME_BITS'd1741371327, `RNS_PRIME_BITS'd1691402272},
			'{`RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd411626274, `RNS_PRIME_BITS'd947299019, `RNS_PRIME_BITS'd922955371, `RNS_PRIME_BITS'd717008281, `RNS_PRIME_BITS'd1830111594, `RNS_PRIME_BITS'd934508094, `RNS_PRIME_BITS'd1421205889, `RNS_PRIME_BITS'd449988104, `RNS_PRIME_BITS'd831748033, `RNS_PRIME_BITS'd1508983539},
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd557538557, `RNS_PRIME_BITS'd403490750, `RNS_PRIME_BITS'd1949898690, `RNS_PRIME_BITS'd673824242, `RNS_PRIME_BITS'd2140456654, `RNS_PRIME_BITS'd1593737565, `RNS_PRIME_BITS'd1112187232, `RNS_PRIME_BITS'd662788483, `RNS_PRIME_BITS'd2062326798, `RNS_PRIME_BITS'd620144669},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1816920898, `RNS_PRIME_BITS'd1094384141, `RNS_PRIME_BITS'd1063616161, `RNS_PRIME_BITS'd177646934, `RNS_PRIME_BITS'd637624846, `RNS_PRIME_BITS'd1034000350, `RNS_PRIME_BITS'd852571262, `RNS_PRIME_BITS'd1123662998, `RNS_PRIME_BITS'd1912514370, `RNS_PRIME_BITS'd670503665},
			'{`RNS_PRIME_BITS'd63, `RNS_PRIME_BITS'd810602857, `RNS_PRIME_BITS'd642107402, `RNS_PRIME_BITS'd501835601, `RNS_PRIME_BITS'd2100152087, `RNS_PRIME_BITS'd1434180654, `RNS_PRIME_BITS'd1473546440, `RNS_PRIME_BITS'd1743054513, `RNS_PRIME_BITS'd1061984730, `RNS_PRIME_BITS'd1279046600, `RNS_PRIME_BITS'd672215837},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd1163688274, `RNS_PRIME_BITS'd1975455806, `RNS_PRIME_BITS'd1738868248, `RNS_PRIME_BITS'd1028163680, `RNS_PRIME_BITS'd1948955802, `RNS_PRIME_BITS'd258261909, `RNS_PRIME_BITS'd62044728, `RNS_PRIME_BITS'd2104716124, `RNS_PRIME_BITS'd835813621, `RNS_PRIME_BITS'd2116158518},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd888549505, `RNS_PRIME_BITS'd408379797, `RNS_PRIME_BITS'd1615714950, `RNS_PRIME_BITS'd335193254, `RNS_PRIME_BITS'd778382437, `RNS_PRIME_BITS'd1404999444, `RNS_PRIME_BITS'd2094919334, `RNS_PRIME_BITS'd1000731411, `RNS_PRIME_BITS'd128514056, `RNS_PRIME_BITS'd1308960976},
			'{`RNS_PRIME_BITS'd63, `RNS_PRIME_BITS'd172802360, `RNS_PRIME_BITS'd1084678325, `RNS_PRIME_BITS'd1426773007, `RNS_PRIME_BITS'd2007192057, `RNS_PRIME_BITS'd1534927494, `RNS_PRIME_BITS'd222234031, `RNS_PRIME_BITS'd1014283952, `RNS_PRIME_BITS'd212408013, `RNS_PRIME_BITS'd1040114333, `RNS_PRIME_BITS'd1959840149},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd2042127020, `RNS_PRIME_BITS'd651195968, `RNS_PRIME_BITS'd584785812, `RNS_PRIME_BITS'd1068763318, `RNS_PRIME_BITS'd25286577, `RNS_PRIME_BITS'd499632345, `RNS_PRIME_BITS'd1201946635, `RNS_PRIME_BITS'd1683948373, `RNS_PRIME_BITS'd1259854149, `RNS_PRIME_BITS'd2027011754},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd1762983961, `RNS_PRIME_BITS'd789211527, `RNS_PRIME_BITS'd526958947, `RNS_PRIME_BITS'd1920112950, `RNS_PRIME_BITS'd1354448624, `RNS_PRIME_BITS'd1238627247, `RNS_PRIME_BITS'd423458879, `RNS_PRIME_BITS'd244123768, `RNS_PRIME_BITS'd190083090, `RNS_PRIME_BITS'd1062535998},
			'{`RNS_PRIME_BITS'd108, `RNS_PRIME_BITS'd717204368, `RNS_PRIME_BITS'd1740153951, `RNS_PRIME_BITS'd2053675152, `RNS_PRIME_BITS'd1619873957, `RNS_PRIME_BITS'd1098557552, `RNS_PRIME_BITS'd293082939, `RNS_PRIME_BITS'd960106005, `RNS_PRIME_BITS'd2069633253, `RNS_PRIME_BITS'd1791303388, `RNS_PRIME_BITS'd1447596142},
			'{`RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd442414040, `RNS_PRIME_BITS'd861656642, `RNS_PRIME_BITS'd2072002555, `RNS_PRIME_BITS'd495518099, `RNS_PRIME_BITS'd1540685654, `RNS_PRIME_BITS'd252094518, `RNS_PRIME_BITS'd2028645591, `RNS_PRIME_BITS'd454101729, `RNS_PRIME_BITS'd548035466, `RNS_PRIME_BITS'd633102971},
			'{`RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd1515586327, `RNS_PRIME_BITS'd209328431, `RNS_PRIME_BITS'd199062626, `RNS_PRIME_BITS'd216501055, `RNS_PRIME_BITS'd1067851881, `RNS_PRIME_BITS'd978630716, `RNS_PRIME_BITS'd810337562, `RNS_PRIME_BITS'd349316834, `RNS_PRIME_BITS'd2028063606, `RNS_PRIME_BITS'd1977631120},
			'{`RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd673584767, `RNS_PRIME_BITS'd2093518202, `RNS_PRIME_BITS'd515850055, `RNS_PRIME_BITS'd2131044671, `RNS_PRIME_BITS'd1522324298, `RNS_PRIME_BITS'd977147766, `RNS_PRIME_BITS'd703005940, `RNS_PRIME_BITS'd740167003, `RNS_PRIME_BITS'd2093175003, `RNS_PRIME_BITS'd946997638},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1389424887, `RNS_PRIME_BITS'd1274242658, `RNS_PRIME_BITS'd840113875, `RNS_PRIME_BITS'd1063624443, `RNS_PRIME_BITS'd1102029110, `RNS_PRIME_BITS'd1685500365, `RNS_PRIME_BITS'd1316169586, `RNS_PRIME_BITS'd1874167445, `RNS_PRIME_BITS'd1704965031, `RNS_PRIME_BITS'd64607735},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd1655791428, `RNS_PRIME_BITS'd1159247602, `RNS_PRIME_BITS'd331710730, `RNS_PRIME_BITS'd913810118, `RNS_PRIME_BITS'd539900470, `RNS_PRIME_BITS'd1740981319, `RNS_PRIME_BITS'd1251325324, `RNS_PRIME_BITS'd755696250, `RNS_PRIME_BITS'd827024774, `RNS_PRIME_BITS'd78686657},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd2088195049, `RNS_PRIME_BITS'd708665714, `RNS_PRIME_BITS'd775223620, `RNS_PRIME_BITS'd314320395, `RNS_PRIME_BITS'd147826306, `RNS_PRIME_BITS'd971719585, `RNS_PRIME_BITS'd2063288752, `RNS_PRIME_BITS'd143342128, `RNS_PRIME_BITS'd656153075, `RNS_PRIME_BITS'd1907587086},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1226652846, `RNS_PRIME_BITS'd865333171, `RNS_PRIME_BITS'd17323864, `RNS_PRIME_BITS'd938625563, `RNS_PRIME_BITS'd1295360322, `RNS_PRIME_BITS'd737360518, `RNS_PRIME_BITS'd327518919, `RNS_PRIME_BITS'd1126059694, `RNS_PRIME_BITS'd211407430, `RNS_PRIME_BITS'd1242644929},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd827657271, `RNS_PRIME_BITS'd876119702, `RNS_PRIME_BITS'd740442358, `RNS_PRIME_BITS'd1044814163, `RNS_PRIME_BITS'd1741004815, `RNS_PRIME_BITS'd628729294, `RNS_PRIME_BITS'd45107064, `RNS_PRIME_BITS'd700450461, `RNS_PRIME_BITS'd807147154, `RNS_PRIME_BITS'd2100412248},
			'{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd116243023, `RNS_PRIME_BITS'd233525114, `RNS_PRIME_BITS'd1323042428, `RNS_PRIME_BITS'd221853300, `RNS_PRIME_BITS'd1063263008, `RNS_PRIME_BITS'd1430397227, `RNS_PRIME_BITS'd612303232, `RNS_PRIME_BITS'd414907045, `RNS_PRIME_BITS'd1793464219, `RNS_PRIME_BITS'd1181884623},
			'{`RNS_PRIME_BITS'd204, `RNS_PRIME_BITS'd1125361005, `RNS_PRIME_BITS'd778542540, `RNS_PRIME_BITS'd1825879191, `RNS_PRIME_BITS'd1320621908, `RNS_PRIME_BITS'd571264056, `RNS_PRIME_BITS'd1750534173, `RNS_PRIME_BITS'd904001111, `RNS_PRIME_BITS'd1237892712, `RNS_PRIME_BITS'd1001030037, `RNS_PRIME_BITS'd226656206},
			'{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd37399989, `RNS_PRIME_BITS'd909904965, `RNS_PRIME_BITS'd832520370, `RNS_PRIME_BITS'd1082666971, `RNS_PRIME_BITS'd414110457, `RNS_PRIME_BITS'd1324824695, `RNS_PRIME_BITS'd974950528, `RNS_PRIME_BITS'd739262197, `RNS_PRIME_BITS'd1807779309, `RNS_PRIME_BITS'd1195940513},
			'{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd182718135, `RNS_PRIME_BITS'd1152435134, `RNS_PRIME_BITS'd1421898968, `RNS_PRIME_BITS'd87950801, `RNS_PRIME_BITS'd468197900, `RNS_PRIME_BITS'd59999510, `RNS_PRIME_BITS'd1271929291, `RNS_PRIME_BITS'd1651773790, `RNS_PRIME_BITS'd145339822, `RNS_PRIME_BITS'd355349572},
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd1350809504, `RNS_PRIME_BITS'd802677379, `RNS_PRIME_BITS'd527818842, `RNS_PRIME_BITS'd906622453, `RNS_PRIME_BITS'd1891955955, `RNS_PRIME_BITS'd1881225418, `RNS_PRIME_BITS'd1626737960, `RNS_PRIME_BITS'd1409740065, `RNS_PRIME_BITS'd1392544884, `RNS_PRIME_BITS'd232748340},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd1481600591, `RNS_PRIME_BITS'd197384772, `RNS_PRIME_BITS'd763042000, `RNS_PRIME_BITS'd357978036, `RNS_PRIME_BITS'd1267901905, `RNS_PRIME_BITS'd1581791892, `RNS_PRIME_BITS'd1240265033, `RNS_PRIME_BITS'd445749290, `RNS_PRIME_BITS'd1696450644, `RNS_PRIME_BITS'd128501568},
			'{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd1797772693, `RNS_PRIME_BITS'd331924767, `RNS_PRIME_BITS'd362173682, `RNS_PRIME_BITS'd27368257, `RNS_PRIME_BITS'd594576380, `RNS_PRIME_BITS'd689176117, `RNS_PRIME_BITS'd361974584, `RNS_PRIME_BITS'd740370380, `RNS_PRIME_BITS'd88511865, `RNS_PRIME_BITS'd1108967642},
			'{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd924677876, `RNS_PRIME_BITS'd654623074, `RNS_PRIME_BITS'd85744617, `RNS_PRIME_BITS'd88731529, `RNS_PRIME_BITS'd1042983153, `RNS_PRIME_BITS'd272334075, `RNS_PRIME_BITS'd1003642840, `RNS_PRIME_BITS'd389864086, `RNS_PRIME_BITS'd1408123962, `RNS_PRIME_BITS'd1047500929},
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd166515930, `RNS_PRIME_BITS'd1944916265, `RNS_PRIME_BITS'd276883350, `RNS_PRIME_BITS'd781010873, `RNS_PRIME_BITS'd959141786, `RNS_PRIME_BITS'd578905400, `RNS_PRIME_BITS'd1764453123, `RNS_PRIME_BITS'd1346272431, `RNS_PRIME_BITS'd1785834928, `RNS_PRIME_BITS'd1204949889},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1792308921, `RNS_PRIME_BITS'd2091131312, `RNS_PRIME_BITS'd522632911, `RNS_PRIME_BITS'd1961335097, `RNS_PRIME_BITS'd584344325, `RNS_PRIME_BITS'd376976427, `RNS_PRIME_BITS'd1822873521, `RNS_PRIME_BITS'd1550923118, `RNS_PRIME_BITS'd232419326, `RNS_PRIME_BITS'd1770869656},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd1879712196, `RNS_PRIME_BITS'd1822702762, `RNS_PRIME_BITS'd1919753088, `RNS_PRIME_BITS'd641835156, `RNS_PRIME_BITS'd1643743751, `RNS_PRIME_BITS'd1077448430, `RNS_PRIME_BITS'd26300314, `RNS_PRIME_BITS'd167303702, `RNS_PRIME_BITS'd245375118, `RNS_PRIME_BITS'd327877411},
			'{`RNS_PRIME_BITS'd170, `RNS_PRIME_BITS'd1623030566, `RNS_PRIME_BITS'd1451408470, `RNS_PRIME_BITS'd389144076, `RNS_PRIME_BITS'd515460666, `RNS_PRIME_BITS'd34483084, `RNS_PRIME_BITS'd688152997, `RNS_PRIME_BITS'd1355495851, `RNS_PRIME_BITS'd1577667674, `RNS_PRIME_BITS'd613227965, `RNS_PRIME_BITS'd1369071893},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1589361954, `RNS_PRIME_BITS'd1001988187, `RNS_PRIME_BITS'd874576670, `RNS_PRIME_BITS'd751132843, `RNS_PRIME_BITS'd1333733331, `RNS_PRIME_BITS'd1216464028, `RNS_PRIME_BITS'd604222924, `RNS_PRIME_BITS'd2095261758, `RNS_PRIME_BITS'd1908544630, `RNS_PRIME_BITS'd1188699792},
			'{`RNS_PRIME_BITS'd142, `RNS_PRIME_BITS'd1933927994, `RNS_PRIME_BITS'd96828190, `RNS_PRIME_BITS'd563422019, `RNS_PRIME_BITS'd974215543, `RNS_PRIME_BITS'd860411096, `RNS_PRIME_BITS'd507519969, `RNS_PRIME_BITS'd166651087, `RNS_PRIME_BITS'd2093869483, `RNS_PRIME_BITS'd1025333640, `RNS_PRIME_BITS'd1199382415},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd397643835, `RNS_PRIME_BITS'd1685579513, `RNS_PRIME_BITS'd1666264534, `RNS_PRIME_BITS'd2144701602, `RNS_PRIME_BITS'd487899691, `RNS_PRIME_BITS'd1344231914, `RNS_PRIME_BITS'd2133536225, `RNS_PRIME_BITS'd1797143825, `RNS_PRIME_BITS'd1967768157, `RNS_PRIME_BITS'd60717247},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd2010011810, `RNS_PRIME_BITS'd1196526663, `RNS_PRIME_BITS'd884777343, `RNS_PRIME_BITS'd895985273, `RNS_PRIME_BITS'd121857223, `RNS_PRIME_BITS'd1757270257, `RNS_PRIME_BITS'd2015454239, `RNS_PRIME_BITS'd1170375999, `RNS_PRIME_BITS'd1902435066, `RNS_PRIME_BITS'd681760182},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd1612149840, `RNS_PRIME_BITS'd477872052, `RNS_PRIME_BITS'd1697400104, `RNS_PRIME_BITS'd1180251613, `RNS_PRIME_BITS'd841422337, `RNS_PRIME_BITS'd1023332073, `RNS_PRIME_BITS'd1053301351, `RNS_PRIME_BITS'd1129973989, `RNS_PRIME_BITS'd305632012, `RNS_PRIME_BITS'd1180561195},
			'{`RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd684810114, `RNS_PRIME_BITS'd159616922, `RNS_PRIME_BITS'd1123921359, `RNS_PRIME_BITS'd1131293257, `RNS_PRIME_BITS'd588800603, `RNS_PRIME_BITS'd925273517, `RNS_PRIME_BITS'd357125827, `RNS_PRIME_BITS'd2053889957, `RNS_PRIME_BITS'd1396416986, `RNS_PRIME_BITS'd1102749471},
			'{`RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd777815011, `RNS_PRIME_BITS'd1633536392, `RNS_PRIME_BITS'd200207179, `RNS_PRIME_BITS'd880121864, `RNS_PRIME_BITS'd1128690021, `RNS_PRIME_BITS'd187488433, `RNS_PRIME_BITS'd1066979046, `RNS_PRIME_BITS'd261956602, `RNS_PRIME_BITS'd766165801, `RNS_PRIME_BITS'd1276067568},
			'{`RNS_PRIME_BITS'd148, `RNS_PRIME_BITS'd1012466243, `RNS_PRIME_BITS'd966034172, `RNS_PRIME_BITS'd139496663, `RNS_PRIME_BITS'd473551751, `RNS_PRIME_BITS'd250893963, `RNS_PRIME_BITS'd746649673, `RNS_PRIME_BITS'd360747560, `RNS_PRIME_BITS'd1477540983, `RNS_PRIME_BITS'd268428551, `RNS_PRIME_BITS'd1274955083}
		},
		'{
			'{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd121221212, `RNS_PRIME_BITS'd1951255688, `RNS_PRIME_BITS'd1301379771, `RNS_PRIME_BITS'd475722016, `RNS_PRIME_BITS'd1304943171, `RNS_PRIME_BITS'd2022962164, `RNS_PRIME_BITS'd1560324161, `RNS_PRIME_BITS'd495684847, `RNS_PRIME_BITS'd1336604873, `RNS_PRIME_BITS'd1416054658},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd1601576126, `RNS_PRIME_BITS'd1069627163, `RNS_PRIME_BITS'd791263671, `RNS_PRIME_BITS'd1452976862, `RNS_PRIME_BITS'd1140310033, `RNS_PRIME_BITS'd790719143, `RNS_PRIME_BITS'd62744675, `RNS_PRIME_BITS'd233100956, `RNS_PRIME_BITS'd899412076, `RNS_PRIME_BITS'd729684010},
			'{`RNS_PRIME_BITS'd65, `RNS_PRIME_BITS'd326679050, `RNS_PRIME_BITS'd968300213, `RNS_PRIME_BITS'd347546755, `RNS_PRIME_BITS'd1185034959, `RNS_PRIME_BITS'd766182269, `RNS_PRIME_BITS'd703271330, `RNS_PRIME_BITS'd2043951564, `RNS_PRIME_BITS'd1844685748, `RNS_PRIME_BITS'd992110879, `RNS_PRIME_BITS'd973336482},
			'{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd1655970335, `RNS_PRIME_BITS'd2129215425, `RNS_PRIME_BITS'd194179222, `RNS_PRIME_BITS'd725198308, `RNS_PRIME_BITS'd1690125207, `RNS_PRIME_BITS'd1439141073, `RNS_PRIME_BITS'd829492529, `RNS_PRIME_BITS'd737320529, `RNS_PRIME_BITS'd255735728, `RNS_PRIME_BITS'd684386041},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd157062667, `RNS_PRIME_BITS'd2014579820, `RNS_PRIME_BITS'd720613023, `RNS_PRIME_BITS'd1489131268, `RNS_PRIME_BITS'd296553590, `RNS_PRIME_BITS'd1126465511, `RNS_PRIME_BITS'd1320190940, `RNS_PRIME_BITS'd578790694, `RNS_PRIME_BITS'd805023131, `RNS_PRIME_BITS'd1859743606},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd1512730238, `RNS_PRIME_BITS'd1718983884, `RNS_PRIME_BITS'd932187246, `RNS_PRIME_BITS'd546661568, `RNS_PRIME_BITS'd784683520, `RNS_PRIME_BITS'd1477725496, `RNS_PRIME_BITS'd1919984576, `RNS_PRIME_BITS'd1890061370, `RNS_PRIME_BITS'd1597149649, `RNS_PRIME_BITS'd2024875218},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd58767579, `RNS_PRIME_BITS'd183578801, `RNS_PRIME_BITS'd725278730, `RNS_PRIME_BITS'd817057599, `RNS_PRIME_BITS'd694543133, `RNS_PRIME_BITS'd169880457, `RNS_PRIME_BITS'd173779742, `RNS_PRIME_BITS'd796141820, `RNS_PRIME_BITS'd1537592220, `RNS_PRIME_BITS'd1543620201},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1934703216, `RNS_PRIME_BITS'd112323919, `RNS_PRIME_BITS'd129495794, `RNS_PRIME_BITS'd931408875, `RNS_PRIME_BITS'd1959738602, `RNS_PRIME_BITS'd926821812, `RNS_PRIME_BITS'd1793200784, `RNS_PRIME_BITS'd1707534163, `RNS_PRIME_BITS'd1896505479, `RNS_PRIME_BITS'd1312281082},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd1565551690, `RNS_PRIME_BITS'd1234193164, `RNS_PRIME_BITS'd802150725, `RNS_PRIME_BITS'd483390414, `RNS_PRIME_BITS'd1964626658, `RNS_PRIME_BITS'd1513234015, `RNS_PRIME_BITS'd2055597025, `RNS_PRIME_BITS'd1730285342, `RNS_PRIME_BITS'd1609634173, `RNS_PRIME_BITS'd1714344332},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd410571370, `RNS_PRIME_BITS'd305318676, `RNS_PRIME_BITS'd921460341, `RNS_PRIME_BITS'd1563432877, `RNS_PRIME_BITS'd1824202795, `RNS_PRIME_BITS'd1724154053, `RNS_PRIME_BITS'd562881691, `RNS_PRIME_BITS'd291376216, `RNS_PRIME_BITS'd381284298, `RNS_PRIME_BITS'd2133100130},
			'{`RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd185532521, `RNS_PRIME_BITS'd210377531, `RNS_PRIME_BITS'd1088514056, `RNS_PRIME_BITS'd1207593828, `RNS_PRIME_BITS'd1368276642, `RNS_PRIME_BITS'd1755245263, `RNS_PRIME_BITS'd1505356531, `RNS_PRIME_BITS'd1784191888, `RNS_PRIME_BITS'd2063241513, `RNS_PRIME_BITS'd1503529633},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd2009319159, `RNS_PRIME_BITS'd1229919801, `RNS_PRIME_BITS'd1795945488, `RNS_PRIME_BITS'd85716195, `RNS_PRIME_BITS'd1566477027, `RNS_PRIME_BITS'd911632031, `RNS_PRIME_BITS'd2135572978, `RNS_PRIME_BITS'd73561723, `RNS_PRIME_BITS'd782234307, `RNS_PRIME_BITS'd62625341},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd1784889968, `RNS_PRIME_BITS'd841743165, `RNS_PRIME_BITS'd217321653, `RNS_PRIME_BITS'd288776839, `RNS_PRIME_BITS'd134132771, `RNS_PRIME_BITS'd749432266, `RNS_PRIME_BITS'd979855439, `RNS_PRIME_BITS'd1009168827, `RNS_PRIME_BITS'd316129983, `RNS_PRIME_BITS'd1490819683},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd69000838, `RNS_PRIME_BITS'd1105019986, `RNS_PRIME_BITS'd1605397288, `RNS_PRIME_BITS'd988803610, `RNS_PRIME_BITS'd2032579412, `RNS_PRIME_BITS'd1332347564, `RNS_PRIME_BITS'd1727567918, `RNS_PRIME_BITS'd283208212, `RNS_PRIME_BITS'd1521763375, `RNS_PRIME_BITS'd72615413},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1850735661, `RNS_PRIME_BITS'd1178071244, `RNS_PRIME_BITS'd1220215830, `RNS_PRIME_BITS'd1534880030, `RNS_PRIME_BITS'd733482146, `RNS_PRIME_BITS'd974234921, `RNS_PRIME_BITS'd197915233, `RNS_PRIME_BITS'd2114199393, `RNS_PRIME_BITS'd1360097077, `RNS_PRIME_BITS'd838270822},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd724286314, `RNS_PRIME_BITS'd2003201690, `RNS_PRIME_BITS'd207962778, `RNS_PRIME_BITS'd479127032, `RNS_PRIME_BITS'd448895285, `RNS_PRIME_BITS'd1795131171, `RNS_PRIME_BITS'd327135205, `RNS_PRIME_BITS'd12943876, `RNS_PRIME_BITS'd791403803, `RNS_PRIME_BITS'd11758094},
			'{`RNS_PRIME_BITS'd5, `RNS_PRIME_BITS'd1718979089, `RNS_PRIME_BITS'd615502449, `RNS_PRIME_BITS'd1481194129, `RNS_PRIME_BITS'd1052637578, `RNS_PRIME_BITS'd560954237, `RNS_PRIME_BITS'd1512751646, `RNS_PRIME_BITS'd2146798395, `RNS_PRIME_BITS'd1416251710, `RNS_PRIME_BITS'd1872662830, `RNS_PRIME_BITS'd1463295855},
			'{`RNS_PRIME_BITS'd171, `RNS_PRIME_BITS'd308885162, `RNS_PRIME_BITS'd243444592, `RNS_PRIME_BITS'd497472652, `RNS_PRIME_BITS'd1004743023, `RNS_PRIME_BITS'd1735683645, `RNS_PRIME_BITS'd1884229621, `RNS_PRIME_BITS'd608637773, `RNS_PRIME_BITS'd273321707, `RNS_PRIME_BITS'd196921081, `RNS_PRIME_BITS'd571284636},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd1887349786, `RNS_PRIME_BITS'd1780505790, `RNS_PRIME_BITS'd436633042, `RNS_PRIME_BITS'd1025292879, `RNS_PRIME_BITS'd217614169, `RNS_PRIME_BITS'd2126325213, `RNS_PRIME_BITS'd1536440905, `RNS_PRIME_BITS'd1397065393, `RNS_PRIME_BITS'd452711235, `RNS_PRIME_BITS'd440954482},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd34776507, `RNS_PRIME_BITS'd1879283380, `RNS_PRIME_BITS'd22898680, `RNS_PRIME_BITS'd889843268, `RNS_PRIME_BITS'd1221747482, `RNS_PRIME_BITS'd1392452286, `RNS_PRIME_BITS'd141645892, `RNS_PRIME_BITS'd88708159, `RNS_PRIME_BITS'd1116579621, `RNS_PRIME_BITS'd1953952519},
			'{`RNS_PRIME_BITS'd126, `RNS_PRIME_BITS'd156492078, `RNS_PRIME_BITS'd270815508, `RNS_PRIME_BITS'd24008909, `RNS_PRIME_BITS'd619028259, `RNS_PRIME_BITS'd1310197468, `RNS_PRIME_BITS'd1462189361, `RNS_PRIME_BITS'd357736511, `RNS_PRIME_BITS'd427467901, `RNS_PRIME_BITS'd1575952606, `RNS_PRIME_BITS'd1003128530},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd14351213, `RNS_PRIME_BITS'd1253972066, `RNS_PRIME_BITS'd414934004, `RNS_PRIME_BITS'd1608707256, `RNS_PRIME_BITS'd134115981, `RNS_PRIME_BITS'd355052224, `RNS_PRIME_BITS'd283938992, `RNS_PRIME_BITS'd1329188123, `RNS_PRIME_BITS'd38360962, `RNS_PRIME_BITS'd1645607187},
			'{`RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd412298267, `RNS_PRIME_BITS'd65261823, `RNS_PRIME_BITS'd1100206669, `RNS_PRIME_BITS'd603850546, `RNS_PRIME_BITS'd709106040, `RNS_PRIME_BITS'd935575719, `RNS_PRIME_BITS'd1316593946, `RNS_PRIME_BITS'd1941035192, `RNS_PRIME_BITS'd551493654, `RNS_PRIME_BITS'd1744002825},
			'{`RNS_PRIME_BITS'd65, `RNS_PRIME_BITS'd303890218, `RNS_PRIME_BITS'd1613003273, `RNS_PRIME_BITS'd540284217, `RNS_PRIME_BITS'd574403678, `RNS_PRIME_BITS'd529231709, `RNS_PRIME_BITS'd484741481, `RNS_PRIME_BITS'd1615463718, `RNS_PRIME_BITS'd672420762, `RNS_PRIME_BITS'd1599202786, `RNS_PRIME_BITS'd1071684640},
			'{`RNS_PRIME_BITS'd20, `RNS_PRIME_BITS'd1775450753, `RNS_PRIME_BITS'd1857112608, `RNS_PRIME_BITS'd1617605667, `RNS_PRIME_BITS'd1839976754, `RNS_PRIME_BITS'd43053002, `RNS_PRIME_BITS'd656193025, `RNS_PRIME_BITS'd218081952, `RNS_PRIME_BITS'd676941754, `RNS_PRIME_BITS'd1513263976, `RNS_PRIME_BITS'd2001171338},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd670458327, `RNS_PRIME_BITS'd474780789, `RNS_PRIME_BITS'd2087852772, `RNS_PRIME_BITS'd41671733, `RNS_PRIME_BITS'd1622132522, `RNS_PRIME_BITS'd1609915920, `RNS_PRIME_BITS'd1336368087, `RNS_PRIME_BITS'd464767730, `RNS_PRIME_BITS'd832926815, `RNS_PRIME_BITS'd1379050699},
			'{`RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd1122412345, `RNS_PRIME_BITS'd1869302691, `RNS_PRIME_BITS'd1779206133, `RNS_PRIME_BITS'd2062985667, `RNS_PRIME_BITS'd369476668, `RNS_PRIME_BITS'd2091749166, `RNS_PRIME_BITS'd1038074180, `RNS_PRIME_BITS'd1950443775, `RNS_PRIME_BITS'd240106665, `RNS_PRIME_BITS'd1766951167},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd613024489, `RNS_PRIME_BITS'd1129781523, `RNS_PRIME_BITS'd1666167746, `RNS_PRIME_BITS'd327213962, `RNS_PRIME_BITS'd1190746592, `RNS_PRIME_BITS'd850567895, `RNS_PRIME_BITS'd1692714702, `RNS_PRIME_BITS'd1148099677, `RNS_PRIME_BITS'd1449950455, `RNS_PRIME_BITS'd502961038},
			'{`RNS_PRIME_BITS'd240, `RNS_PRIME_BITS'd461719806, `RNS_PRIME_BITS'd1769354757, `RNS_PRIME_BITS'd894704121, `RNS_PRIME_BITS'd2036967849, `RNS_PRIME_BITS'd101539305, `RNS_PRIME_BITS'd1560357209, `RNS_PRIME_BITS'd1901066514, `RNS_PRIME_BITS'd193016899, `RNS_PRIME_BITS'd1185201792, `RNS_PRIME_BITS'd810800789},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd1781990923, `RNS_PRIME_BITS'd952845231, `RNS_PRIME_BITS'd917663953, `RNS_PRIME_BITS'd20261753, `RNS_PRIME_BITS'd1658234054, `RNS_PRIME_BITS'd598108465, `RNS_PRIME_BITS'd429826561, `RNS_PRIME_BITS'd337240893, `RNS_PRIME_BITS'd1625038773, `RNS_PRIME_BITS'd1719477231},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd1051970377, `RNS_PRIME_BITS'd766984126, `RNS_PRIME_BITS'd298498072, `RNS_PRIME_BITS'd606643384, `RNS_PRIME_BITS'd1447967229, `RNS_PRIME_BITS'd1176830711, `RNS_PRIME_BITS'd742410082, `RNS_PRIME_BITS'd1452847844, `RNS_PRIME_BITS'd360669530, `RNS_PRIME_BITS'd2063959897},
			'{`RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd1101984053, `RNS_PRIME_BITS'd2056771642, `RNS_PRIME_BITS'd1988938968, `RNS_PRIME_BITS'd944305037, `RNS_PRIME_BITS'd1330832185, `RNS_PRIME_BITS'd1422542589, `RNS_PRIME_BITS'd1702452074, `RNS_PRIME_BITS'd693519816, `RNS_PRIME_BITS'd1636569039, `RNS_PRIME_BITS'd385451156},
			'{`RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd522300364, `RNS_PRIME_BITS'd785888962, `RNS_PRIME_BITS'd1897585472, `RNS_PRIME_BITS'd960210142, `RNS_PRIME_BITS'd1986820352, `RNS_PRIME_BITS'd288649031, `RNS_PRIME_BITS'd393792544, `RNS_PRIME_BITS'd1434623371, `RNS_PRIME_BITS'd944607389, `RNS_PRIME_BITS'd1271299749},
			'{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd766366547, `RNS_PRIME_BITS'd1247127502, `RNS_PRIME_BITS'd186185856, `RNS_PRIME_BITS'd1409069545, `RNS_PRIME_BITS'd343937695, `RNS_PRIME_BITS'd1618794645, `RNS_PRIME_BITS'd484565289, `RNS_PRIME_BITS'd135888231, `RNS_PRIME_BITS'd997014915, `RNS_PRIME_BITS'd2048649959},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1275607494, `RNS_PRIME_BITS'd279296353, `RNS_PRIME_BITS'd621264063, `RNS_PRIME_BITS'd377104429, `RNS_PRIME_BITS'd165204523, `RNS_PRIME_BITS'd1508749193, `RNS_PRIME_BITS'd1000657425, `RNS_PRIME_BITS'd891529147, `RNS_PRIME_BITS'd1362879603, `RNS_PRIME_BITS'd2104333727},
			'{`RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd366663080, `RNS_PRIME_BITS'd1618498371, `RNS_PRIME_BITS'd319379119, `RNS_PRIME_BITS'd1065749455, `RNS_PRIME_BITS'd1802523180, `RNS_PRIME_BITS'd1629327637, `RNS_PRIME_BITS'd536813181, `RNS_PRIME_BITS'd2033954784, `RNS_PRIME_BITS'd1419510241, `RNS_PRIME_BITS'd1233439632},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1917285606, `RNS_PRIME_BITS'd1354469122, `RNS_PRIME_BITS'd370772680, `RNS_PRIME_BITS'd1189173244, `RNS_PRIME_BITS'd821356621, `RNS_PRIME_BITS'd1612690931, `RNS_PRIME_BITS'd1097119822, `RNS_PRIME_BITS'd115562925, `RNS_PRIME_BITS'd980236081, `RNS_PRIME_BITS'd1260705325},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1142067223, `RNS_PRIME_BITS'd887765108, `RNS_PRIME_BITS'd1575195784, `RNS_PRIME_BITS'd1566828770, `RNS_PRIME_BITS'd964806824, `RNS_PRIME_BITS'd1350156916, `RNS_PRIME_BITS'd578019889, `RNS_PRIME_BITS'd1384217071, `RNS_PRIME_BITS'd1438278851, `RNS_PRIME_BITS'd1247488765},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1612288038, `RNS_PRIME_BITS'd478496983, `RNS_PRIME_BITS'd1839123021, `RNS_PRIME_BITS'd34067692, `RNS_PRIME_BITS'd1732287927, `RNS_PRIME_BITS'd1909307538, `RNS_PRIME_BITS'd2065185447, `RNS_PRIME_BITS'd897247067, `RNS_PRIME_BITS'd1359706325, `RNS_PRIME_BITS'd1081432982},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd1413194767, `RNS_PRIME_BITS'd401082621, `RNS_PRIME_BITS'd995710083, `RNS_PRIME_BITS'd2036702364, `RNS_PRIME_BITS'd691438769, `RNS_PRIME_BITS'd1491012800, `RNS_PRIME_BITS'd586190011, `RNS_PRIME_BITS'd553405390, `RNS_PRIME_BITS'd241445354, `RNS_PRIME_BITS'd1518161160},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd860850265, `RNS_PRIME_BITS'd1632694784, `RNS_PRIME_BITS'd2138508508, `RNS_PRIME_BITS'd1465058960, `RNS_PRIME_BITS'd829723164, `RNS_PRIME_BITS'd1466257475, `RNS_PRIME_BITS'd611819455, `RNS_PRIME_BITS'd1167998434, `RNS_PRIME_BITS'd631094293, `RNS_PRIME_BITS'd1824186488},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd691990357, `RNS_PRIME_BITS'd1871602326, `RNS_PRIME_BITS'd1253902905, `RNS_PRIME_BITS'd1515478300, `RNS_PRIME_BITS'd1238819032, `RNS_PRIME_BITS'd360154198, `RNS_PRIME_BITS'd1093198667, `RNS_PRIME_BITS'd999911929, `RNS_PRIME_BITS'd706404180, `RNS_PRIME_BITS'd516355116},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd1707748512, `RNS_PRIME_BITS'd1685391667, `RNS_PRIME_BITS'd1698637754, `RNS_PRIME_BITS'd191781474, `RNS_PRIME_BITS'd1497369485, `RNS_PRIME_BITS'd1285710995, `RNS_PRIME_BITS'd743889193, `RNS_PRIME_BITS'd1584878257, `RNS_PRIME_BITS'd647867191, `RNS_PRIME_BITS'd185077071},
			'{`RNS_PRIME_BITS'd76, `RNS_PRIME_BITS'd921242189, `RNS_PRIME_BITS'd657401959, `RNS_PRIME_BITS'd2113054314, `RNS_PRIME_BITS'd97598861, `RNS_PRIME_BITS'd2008697854, `RNS_PRIME_BITS'd527524065, `RNS_PRIME_BITS'd531938748, `RNS_PRIME_BITS'd1185099191, `RNS_PRIME_BITS'd1566650882, `RNS_PRIME_BITS'd1058810141},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd1242612921, `RNS_PRIME_BITS'd166050149, `RNS_PRIME_BITS'd1458366391, `RNS_PRIME_BITS'd1677518012, `RNS_PRIME_BITS'd1467911807, `RNS_PRIME_BITS'd1915522038, `RNS_PRIME_BITS'd1459482010, `RNS_PRIME_BITS'd1446917857, `RNS_PRIME_BITS'd1748614482, `RNS_PRIME_BITS'd1362061942},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd302446774, `RNS_PRIME_BITS'd58933664, `RNS_PRIME_BITS'd489650786, `RNS_PRIME_BITS'd1983885555, `RNS_PRIME_BITS'd318807824, `RNS_PRIME_BITS'd953014828, `RNS_PRIME_BITS'd1046493451, `RNS_PRIME_BITS'd2086293796, `RNS_PRIME_BITS'd780343976, `RNS_PRIME_BITS'd340002060},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd892721966, `RNS_PRIME_BITS'd111645947, `RNS_PRIME_BITS'd1759569081, `RNS_PRIME_BITS'd899965364, `RNS_PRIME_BITS'd307472003, `RNS_PRIME_BITS'd812581241, `RNS_PRIME_BITS'd1598588439, `RNS_PRIME_BITS'd731382113, `RNS_PRIME_BITS'd35554928, `RNS_PRIME_BITS'd1353203382},
			'{`RNS_PRIME_BITS'd14, `RNS_PRIME_BITS'd1853439910, `RNS_PRIME_BITS'd1141473089, `RNS_PRIME_BITS'd1666367350, `RNS_PRIME_BITS'd77511693, `RNS_PRIME_BITS'd855761441, `RNS_PRIME_BITS'd1536620204, `RNS_PRIME_BITS'd8796677, `RNS_PRIME_BITS'd146503383, `RNS_PRIME_BITS'd1824010209, `RNS_PRIME_BITS'd1378324098},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd1582359229, `RNS_PRIME_BITS'd1593121149, `RNS_PRIME_BITS'd2143278437, `RNS_PRIME_BITS'd1013199975, `RNS_PRIME_BITS'd480414426, `RNS_PRIME_BITS'd879934074, `RNS_PRIME_BITS'd1135145037, `RNS_PRIME_BITS'd42734978, `RNS_PRIME_BITS'd888716610, `RNS_PRIME_BITS'd765729092},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd184374192, `RNS_PRIME_BITS'd1537864809, `RNS_PRIME_BITS'd20173061, `RNS_PRIME_BITS'd1313606139, `RNS_PRIME_BITS'd932877088, `RNS_PRIME_BITS'd1460394645, `RNS_PRIME_BITS'd1662115500, `RNS_PRIME_BITS'd446878760, `RNS_PRIME_BITS'd348129187, `RNS_PRIME_BITS'd1280849769},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd1122833377, `RNS_PRIME_BITS'd1870409211, `RNS_PRIME_BITS'd420931038, `RNS_PRIME_BITS'd292120676, `RNS_PRIME_BITS'd1342714626, `RNS_PRIME_BITS'd259174392, `RNS_PRIME_BITS'd1835705299, `RNS_PRIME_BITS'd1248797026, `RNS_PRIME_BITS'd1032633350, `RNS_PRIME_BITS'd1029122214},
			'{`RNS_PRIME_BITS'd163, `RNS_PRIME_BITS'd1389658896, `RNS_PRIME_BITS'd947694778, `RNS_PRIME_BITS'd1894638033, `RNS_PRIME_BITS'd1324860415, `RNS_PRIME_BITS'd1915883999, `RNS_PRIME_BITS'd142088715, `RNS_PRIME_BITS'd165331640, `RNS_PRIME_BITS'd29587290, `RNS_PRIME_BITS'd178714264, `RNS_PRIME_BITS'd1653223470},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd644147692, `RNS_PRIME_BITS'd1035420420, `RNS_PRIME_BITS'd1038371180, `RNS_PRIME_BITS'd1518086210, `RNS_PRIME_BITS'd1127088856, `RNS_PRIME_BITS'd224346910, `RNS_PRIME_BITS'd1504595496, `RNS_PRIME_BITS'd342209808, `RNS_PRIME_BITS'd346406331, `RNS_PRIME_BITS'd1493254837},
			'{`RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd1598820713, `RNS_PRIME_BITS'd901199633, `RNS_PRIME_BITS'd393797718, `RNS_PRIME_BITS'd1338979811, `RNS_PRIME_BITS'd161984477, `RNS_PRIME_BITS'd1896237317, `RNS_PRIME_BITS'd848963471, `RNS_PRIME_BITS'd1959536308, `RNS_PRIME_BITS'd1041623424, `RNS_PRIME_BITS'd845134363},
			'{`RNS_PRIME_BITS'd148, `RNS_PRIME_BITS'd1244121150, `RNS_PRIME_BITS'd955491936, `RNS_PRIME_BITS'd484297377, `RNS_PRIME_BITS'd1608749955, `RNS_PRIME_BITS'd76028533, `RNS_PRIME_BITS'd719142789, `RNS_PRIME_BITS'd965635702, `RNS_PRIME_BITS'd1768579328, `RNS_PRIME_BITS'd1663878682, `RNS_PRIME_BITS'd648275179},
			'{`RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd314669877, `RNS_PRIME_BITS'd1767628276, `RNS_PRIME_BITS'd126651183, `RNS_PRIME_BITS'd1410092720, `RNS_PRIME_BITS'd1631999985, `RNS_PRIME_BITS'd1895397156, `RNS_PRIME_BITS'd1018403627, `RNS_PRIME_BITS'd937053505, `RNS_PRIME_BITS'd1200609512, `RNS_PRIME_BITS'd92628929},
			'{`RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd1779270796, `RNS_PRIME_BITS'd1025291671, `RNS_PRIME_BITS'd1691511185, `RNS_PRIME_BITS'd781019140, `RNS_PRIME_BITS'd1271972833, `RNS_PRIME_BITS'd1592234781, `RNS_PRIME_BITS'd1624205452, `RNS_PRIME_BITS'd1406368702, `RNS_PRIME_BITS'd1268145017, `RNS_PRIME_BITS'd2040373124},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd1032842354, `RNS_PRIME_BITS'd1310312155, `RNS_PRIME_BITS'd1313883967, `RNS_PRIME_BITS'd894266693, `RNS_PRIME_BITS'd1787601205, `RNS_PRIME_BITS'd1269169829, `RNS_PRIME_BITS'd591727438, `RNS_PRIME_BITS'd137692414, `RNS_PRIME_BITS'd1224380143, `RNS_PRIME_BITS'd1703081266},
			'{`RNS_PRIME_BITS'd156, `RNS_PRIME_BITS'd416494418, `RNS_PRIME_BITS'd1626329157, `RNS_PRIME_BITS'd1620368821, `RNS_PRIME_BITS'd1269472365, `RNS_PRIME_BITS'd1068673104, `RNS_PRIME_BITS'd2133688296, `RNS_PRIME_BITS'd570888719, `RNS_PRIME_BITS'd608800642, `RNS_PRIME_BITS'd2060071179, `RNS_PRIME_BITS'd1193510543},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd1637868274, `RNS_PRIME_BITS'd1888034906, `RNS_PRIME_BITS'd213982373, `RNS_PRIME_BITS'd412024193, `RNS_PRIME_BITS'd1439650188, `RNS_PRIME_BITS'd197532198, `RNS_PRIME_BITS'd1588013712, `RNS_PRIME_BITS'd2140570198, `RNS_PRIME_BITS'd1208345422, `RNS_PRIME_BITS'd379831942},
			'{`RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd1409085233, `RNS_PRIME_BITS'd1165606570, `RNS_PRIME_BITS'd1636048528, `RNS_PRIME_BITS'd1746052191, `RNS_PRIME_BITS'd2071151476, `RNS_PRIME_BITS'd683031429, `RNS_PRIME_BITS'd2144523196, `RNS_PRIME_BITS'd435307280, `RNS_PRIME_BITS'd1348723726, `RNS_PRIME_BITS'd1419699817},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd1956759644, `RNS_PRIME_BITS'd1814522908, `RNS_PRIME_BITS'd1987475675, `RNS_PRIME_BITS'd1376594889, `RNS_PRIME_BITS'd1574194848, `RNS_PRIME_BITS'd996378142, `RNS_PRIME_BITS'd619984418, `RNS_PRIME_BITS'd1345021853, `RNS_PRIME_BITS'd25451369, `RNS_PRIME_BITS'd1226304744},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1123921442, `RNS_PRIME_BITS'd133591630, `RNS_PRIME_BITS'd436203089, `RNS_PRIME_BITS'd1021951280, `RNS_PRIME_BITS'd426624464, `RNS_PRIME_BITS'd2137338800, `RNS_PRIME_BITS'd468796009, `RNS_PRIME_BITS'd560685756, `RNS_PRIME_BITS'd758064231, `RNS_PRIME_BITS'd1286624983},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd512825721, `RNS_PRIME_BITS'd901081071, `RNS_PRIME_BITS'd724486466, `RNS_PRIME_BITS'd1661050834, `RNS_PRIME_BITS'd1557532595, `RNS_PRIME_BITS'd649773421, `RNS_PRIME_BITS'd2119956614, `RNS_PRIME_BITS'd405402303, `RNS_PRIME_BITS'd2082990312, `RNS_PRIME_BITS'd956294042}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd206089988, `RNS_PRIME_BITS'd390004685, `RNS_PRIME_BITS'd2133402292, `RNS_PRIME_BITS'd1176399385, `RNS_PRIME_BITS'd27008538, `RNS_PRIME_BITS'd1374772353, `RNS_PRIME_BITS'd593287819, `RNS_PRIME_BITS'd471748892, `RNS_PRIME_BITS'd2009838358, `RNS_PRIME_BITS'd786005650},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1481290386, `RNS_PRIME_BITS'd317099186, `RNS_PRIME_BITS'd338271695, `RNS_PRIME_BITS'd1167722141, `RNS_PRIME_BITS'd2115762618, `RNS_PRIME_BITS'd2008014779, `RNS_PRIME_BITS'd606245044, `RNS_PRIME_BITS'd558567039, `RNS_PRIME_BITS'd127877830, `RNS_PRIME_BITS'd607674041},
			'{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd1127866326, `RNS_PRIME_BITS'd1258939673, `RNS_PRIME_BITS'd1562712308, `RNS_PRIME_BITS'd2144011172, `RNS_PRIME_BITS'd323628270, `RNS_PRIME_BITS'd454518980, `RNS_PRIME_BITS'd701832282, `RNS_PRIME_BITS'd590910916, `RNS_PRIME_BITS'd265866377, `RNS_PRIME_BITS'd84978718},
			'{`RNS_PRIME_BITS'd12, `RNS_PRIME_BITS'd1661390003, `RNS_PRIME_BITS'd965921938, `RNS_PRIME_BITS'd491762016, `RNS_PRIME_BITS'd184943715, `RNS_PRIME_BITS'd1782371355, `RNS_PRIME_BITS'd1746993936, `RNS_PRIME_BITS'd694610233, `RNS_PRIME_BITS'd2015168746, `RNS_PRIME_BITS'd73433080, `RNS_PRIME_BITS'd1036378145},
			'{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd512965494, `RNS_PRIME_BITS'd454617685, `RNS_PRIME_BITS'd1886170279, `RNS_PRIME_BITS'd1430774728, `RNS_PRIME_BITS'd300254645, `RNS_PRIME_BITS'd916609989, `RNS_PRIME_BITS'd885318545, `RNS_PRIME_BITS'd2108738422, `RNS_PRIME_BITS'd15257296, `RNS_PRIME_BITS'd981938093},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd127450082, `RNS_PRIME_BITS'd419116467, `RNS_PRIME_BITS'd613430365, `RNS_PRIME_BITS'd692360395, `RNS_PRIME_BITS'd1784227505, `RNS_PRIME_BITS'd1287280376, `RNS_PRIME_BITS'd1471130847, `RNS_PRIME_BITS'd1268444775, `RNS_PRIME_BITS'd1621336831, `RNS_PRIME_BITS'd161770554},
			'{`RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd2026216472, `RNS_PRIME_BITS'd678712620, `RNS_PRIME_BITS'd574586147, `RNS_PRIME_BITS'd1783737920, `RNS_PRIME_BITS'd812999431, `RNS_PRIME_BITS'd1193916047, `RNS_PRIME_BITS'd931836127, `RNS_PRIME_BITS'd1920769855, `RNS_PRIME_BITS'd1155470089, `RNS_PRIME_BITS'd1361464949},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd1478405719, `RNS_PRIME_BITS'd1043196050, `RNS_PRIME_BITS'd1451416784, `RNS_PRIME_BITS'd583244220, `RNS_PRIME_BITS'd1675854177, `RNS_PRIME_BITS'd2132902663, `RNS_PRIME_BITS'd1812219819, `RNS_PRIME_BITS'd1646962751, `RNS_PRIME_BITS'd1652512611, `RNS_PRIME_BITS'd1018382043},
			'{`RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd138920971, `RNS_PRIME_BITS'd2071963271, `RNS_PRIME_BITS'd1181825851, `RNS_PRIME_BITS'd27424554, `RNS_PRIME_BITS'd2144279937, `RNS_PRIME_BITS'd330725491, `RNS_PRIME_BITS'd1700203170, `RNS_PRIME_BITS'd2026427645, `RNS_PRIME_BITS'd1715103458, `RNS_PRIME_BITS'd184451521},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1846050265, `RNS_PRIME_BITS'd1326479294, `RNS_PRIME_BITS'd790680035, `RNS_PRIME_BITS'd1518767684, `RNS_PRIME_BITS'd897907290, `RNS_PRIME_BITS'd889069269, `RNS_PRIME_BITS'd2001316398, `RNS_PRIME_BITS'd1986237580, `RNS_PRIME_BITS'd2098481783, `RNS_PRIME_BITS'd707282160},
			'{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd27414349, `RNS_PRIME_BITS'd178584342, `RNS_PRIME_BITS'd1078682959, `RNS_PRIME_BITS'd392049398, `RNS_PRIME_BITS'd1599944545, `RNS_PRIME_BITS'd785802467, `RNS_PRIME_BITS'd1282136738, `RNS_PRIME_BITS'd2142001886, `RNS_PRIME_BITS'd1811875993, `RNS_PRIME_BITS'd1840673492},
			'{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd192408700, `RNS_PRIME_BITS'd1814441102, `RNS_PRIME_BITS'd279985613, `RNS_PRIME_BITS'd2054367828, `RNS_PRIME_BITS'd614690586, `RNS_PRIME_BITS'd506236410, `RNS_PRIME_BITS'd1537623707, `RNS_PRIME_BITS'd658932769, `RNS_PRIME_BITS'd1972368337, `RNS_PRIME_BITS'd1595331511},
			'{`RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd1871873258, `RNS_PRIME_BITS'd1784784770, `RNS_PRIME_BITS'd1006656492, `RNS_PRIME_BITS'd1948287082, `RNS_PRIME_BITS'd891824894, `RNS_PRIME_BITS'd265035470, `RNS_PRIME_BITS'd762228546, `RNS_PRIME_BITS'd2084600778, `RNS_PRIME_BITS'd361082005, `RNS_PRIME_BITS'd1856846885},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd1468080625, `RNS_PRIME_BITS'd240616847, `RNS_PRIME_BITS'd2028112262, `RNS_PRIME_BITS'd1842703068, `RNS_PRIME_BITS'd9944733, `RNS_PRIME_BITS'd979107366, `RNS_PRIME_BITS'd490175152, `RNS_PRIME_BITS'd1503350770, `RNS_PRIME_BITS'd949453711, `RNS_PRIME_BITS'd928840176},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd166489078, `RNS_PRIME_BITS'd672096339, `RNS_PRIME_BITS'd315827718, `RNS_PRIME_BITS'd285282683, `RNS_PRIME_BITS'd1731732127, `RNS_PRIME_BITS'd2119893561, `RNS_PRIME_BITS'd88847965, `RNS_PRIME_BITS'd1427275217, `RNS_PRIME_BITS'd1405943937, `RNS_PRIME_BITS'd1490785267},
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd436305949, `RNS_PRIME_BITS'd314734960, `RNS_PRIME_BITS'd810471542, `RNS_PRIME_BITS'd578344224, `RNS_PRIME_BITS'd1191258721, `RNS_PRIME_BITS'd1430639587, `RNS_PRIME_BITS'd1757204757, `RNS_PRIME_BITS'd1766864934, `RNS_PRIME_BITS'd1715573033, `RNS_PRIME_BITS'd310258686},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd68754411, `RNS_PRIME_BITS'd1224190291, `RNS_PRIME_BITS'd789100497, `RNS_PRIME_BITS'd837211010, `RNS_PRIME_BITS'd359037055, `RNS_PRIME_BITS'd2106537032, `RNS_PRIME_BITS'd287847334, `RNS_PRIME_BITS'd1899942205, `RNS_PRIME_BITS'd1868341496, `RNS_PRIME_BITS'd260476724},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd1470870391, `RNS_PRIME_BITS'd234626890, `RNS_PRIME_BITS'd745970360, `RNS_PRIME_BITS'd60566548, `RNS_PRIME_BITS'd859776322, `RNS_PRIME_BITS'd1898770308, `RNS_PRIME_BITS'd1961962090, `RNS_PRIME_BITS'd1741080759, `RNS_PRIME_BITS'd719634577, `RNS_PRIME_BITS'd572099799},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd2016710388, `RNS_PRIME_BITS'd1092936488, `RNS_PRIME_BITS'd1757907351, `RNS_PRIME_BITS'd904206814, `RNS_PRIME_BITS'd1025616058, `RNS_PRIME_BITS'd1073827418, `RNS_PRIME_BITS'd243153673, `RNS_PRIME_BITS'd944881582, `RNS_PRIME_BITS'd2083940145, `RNS_PRIME_BITS'd1258074241},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd581788553, `RNS_PRIME_BITS'd125020229, `RNS_PRIME_BITS'd2076698965, `RNS_PRIME_BITS'd1808305004, `RNS_PRIME_BITS'd455712062, `RNS_PRIME_BITS'd1228612613, `RNS_PRIME_BITS'd1045773729, `RNS_PRIME_BITS'd2008402343, `RNS_PRIME_BITS'd665412424, `RNS_PRIME_BITS'd2118733269},
			'{`RNS_PRIME_BITS'd38, `RNS_PRIME_BITS'd1748485284, `RNS_PRIME_BITS'd1107556707, `RNS_PRIME_BITS'd71501363, `RNS_PRIME_BITS'd1474804469, `RNS_PRIME_BITS'd1670202355, `RNS_PRIME_BITS'd408142158, `RNS_PRIME_BITS'd1890761628, `RNS_PRIME_BITS'd948915769, `RNS_PRIME_BITS'd1287155354, `RNS_PRIME_BITS'd1671739189},
			'{`RNS_PRIME_BITS'd76, `RNS_PRIME_BITS'd1316223137, `RNS_PRIME_BITS'd621618963, `RNS_PRIME_BITS'd1452890027, `RNS_PRIME_BITS'd582927424, `RNS_PRIME_BITS'd657547006, `RNS_PRIME_BITS'd2141310314, `RNS_PRIME_BITS'd1360564711, `RNS_PRIME_BITS'd884515191, `RNS_PRIME_BITS'd2110594296, `RNS_PRIME_BITS'd487216738},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd212712176, `RNS_PRIME_BITS'd1308494355, `RNS_PRIME_BITS'd1919860706, `RNS_PRIME_BITS'd375653914, `RNS_PRIME_BITS'd1291434203, `RNS_PRIME_BITS'd415988957, `RNS_PRIME_BITS'd223806426, `RNS_PRIME_BITS'd779810815, `RNS_PRIME_BITS'd1183003605, `RNS_PRIME_BITS'd2061020856},
			'{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd876273837, `RNS_PRIME_BITS'd1698409806, `RNS_PRIME_BITS'd1760875267, `RNS_PRIME_BITS'd1737143743, `RNS_PRIME_BITS'd1639334704, `RNS_PRIME_BITS'd834681898, `RNS_PRIME_BITS'd1459803520, `RNS_PRIME_BITS'd473080366, `RNS_PRIME_BITS'd260647574, `RNS_PRIME_BITS'd38497828},
			'{`RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd1745546257, `RNS_PRIME_BITS'd110458295, `RNS_PRIME_BITS'd577575810, `RNS_PRIME_BITS'd246195098, `RNS_PRIME_BITS'd342687841, `RNS_PRIME_BITS'd282636999, `RNS_PRIME_BITS'd435438044, `RNS_PRIME_BITS'd1027435600, `RNS_PRIME_BITS'd816939442, `RNS_PRIME_BITS'd1357650647},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd942441668, `RNS_PRIME_BITS'd2137120778, `RNS_PRIME_BITS'd866085588, `RNS_PRIME_BITS'd1186096945, `RNS_PRIME_BITS'd853543971, `RNS_PRIME_BITS'd2030594457, `RNS_PRIME_BITS'd2138514851, `RNS_PRIME_BITS'd2095655488, `RNS_PRIME_BITS'd149947625, `RNS_PRIME_BITS'd1913911692},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd548266251, `RNS_PRIME_BITS'd1470945841, `RNS_PRIME_BITS'd1803569866, `RNS_PRIME_BITS'd1006119583, `RNS_PRIME_BITS'd1547636307, `RNS_PRIME_BITS'd1577553259, `RNS_PRIME_BITS'd607231200, `RNS_PRIME_BITS'd971458844, `RNS_PRIME_BITS'd551260161, `RNS_PRIME_BITS'd149285477},
			'{`RNS_PRIME_BITS'd86, `RNS_PRIME_BITS'd888962987, `RNS_PRIME_BITS'd969284832, `RNS_PRIME_BITS'd89658280, `RNS_PRIME_BITS'd583643777, `RNS_PRIME_BITS'd410243562, `RNS_PRIME_BITS'd346792337, `RNS_PRIME_BITS'd93925565, `RNS_PRIME_BITS'd1315320787, `RNS_PRIME_BITS'd1077545431, `RNS_PRIME_BITS'd1408533358},
			'{`RNS_PRIME_BITS'd85, `RNS_PRIME_BITS'd410514686, `RNS_PRIME_BITS'd147275961, `RNS_PRIME_BITS'd655408583, `RNS_PRIME_BITS'd791763897, `RNS_PRIME_BITS'd687724148, `RNS_PRIME_BITS'd1014515585, `RNS_PRIME_BITS'd727957540, `RNS_PRIME_BITS'd1333568197, `RNS_PRIME_BITS'd964215203, `RNS_PRIME_BITS'd1708346054},
			'{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd1684738999, `RNS_PRIME_BITS'd107265551, `RNS_PRIME_BITS'd308643774, `RNS_PRIME_BITS'd1646796315, `RNS_PRIME_BITS'd1093141154, `RNS_PRIME_BITS'd1235485410, `RNS_PRIME_BITS'd370310755, `RNS_PRIME_BITS'd1275496350, `RNS_PRIME_BITS'd1788816301, `RNS_PRIME_BITS'd735178756},
			'{`RNS_PRIME_BITS'd200, `RNS_PRIME_BITS'd799546255, `RNS_PRIME_BITS'd2071038798, `RNS_PRIME_BITS'd1913639673, `RNS_PRIME_BITS'd268540896, `RNS_PRIME_BITS'd487406235, `RNS_PRIME_BITS'd311170756, `RNS_PRIME_BITS'd1060236694, `RNS_PRIME_BITS'd1822594793, `RNS_PRIME_BITS'd1944803186, `RNS_PRIME_BITS'd179239972},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1818736054, `RNS_PRIME_BITS'd872724654, `RNS_PRIME_BITS'd14711739, `RNS_PRIME_BITS'd304962171, `RNS_PRIME_BITS'd1515823619, `RNS_PRIME_BITS'd2124602952, `RNS_PRIME_BITS'd1656859382, `RNS_PRIME_BITS'd1812906772, `RNS_PRIME_BITS'd1116325779, `RNS_PRIME_BITS'd714902229},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd1166998217, `RNS_PRIME_BITS'd842223466, `RNS_PRIME_BITS'd1258159417, `RNS_PRIME_BITS'd1220543382, `RNS_PRIME_BITS'd1223392789, `RNS_PRIME_BITS'd1073521708, `RNS_PRIME_BITS'd1687185388, `RNS_PRIME_BITS'd2023548152, `RNS_PRIME_BITS'd1469826218, `RNS_PRIME_BITS'd1619805134},
			'{`RNS_PRIME_BITS'd217, `RNS_PRIME_BITS'd1655096059, `RNS_PRIME_BITS'd2073820980, `RNS_PRIME_BITS'd885736280, `RNS_PRIME_BITS'd1870795513, `RNS_PRIME_BITS'd1728535797, `RNS_PRIME_BITS'd666863468, `RNS_PRIME_BITS'd315526539, `RNS_PRIME_BITS'd319594578, `RNS_PRIME_BITS'd2070951595, `RNS_PRIME_BITS'd1617508725},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1782278687, `RNS_PRIME_BITS'd2118156827, `RNS_PRIME_BITS'd1573740365, `RNS_PRIME_BITS'd1615162298, `RNS_PRIME_BITS'd1997859409, `RNS_PRIME_BITS'd1532415036, `RNS_PRIME_BITS'd1240827833, `RNS_PRIME_BITS'd991948942, `RNS_PRIME_BITS'd621853307, `RNS_PRIME_BITS'd1247636363},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd1421696022, `RNS_PRIME_BITS'd2144887985, `RNS_PRIME_BITS'd1420519235, `RNS_PRIME_BITS'd86063047, `RNS_PRIME_BITS'd705404172, `RNS_PRIME_BITS'd722359424, `RNS_PRIME_BITS'd2055553446, `RNS_PRIME_BITS'd2002546155, `RNS_PRIME_BITS'd138407856, `RNS_PRIME_BITS'd2013912438},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd337581797, `RNS_PRIME_BITS'd763318072, `RNS_PRIME_BITS'd899337024, `RNS_PRIME_BITS'd1500078003, `RNS_PRIME_BITS'd1407999938, `RNS_PRIME_BITS'd1790114382, `RNS_PRIME_BITS'd538538241, `RNS_PRIME_BITS'd93762758, `RNS_PRIME_BITS'd1183294065, `RNS_PRIME_BITS'd1533907917},
			'{`RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd1038215496, `RNS_PRIME_BITS'd174334198, `RNS_PRIME_BITS'd1694682842, `RNS_PRIME_BITS'd615955644, `RNS_PRIME_BITS'd171338312, `RNS_PRIME_BITS'd1601406674, `RNS_PRIME_BITS'd1213223166, `RNS_PRIME_BITS'd26879606, `RNS_PRIME_BITS'd154865461, `RNS_PRIME_BITS'd999688025},
			'{`RNS_PRIME_BITS'd15, `RNS_PRIME_BITS'd1285988102, `RNS_PRIME_BITS'd104456546, `RNS_PRIME_BITS'd1487658978, `RNS_PRIME_BITS'd1612781156, `RNS_PRIME_BITS'd1301638207, `RNS_PRIME_BITS'd719273133, `RNS_PRIME_BITS'd774052916, `RNS_PRIME_BITS'd2099739068, `RNS_PRIME_BITS'd1629262359, `RNS_PRIME_BITS'd439444109},
			'{`RNS_PRIME_BITS'd150, `RNS_PRIME_BITS'd1141917621, `RNS_PRIME_BITS'd2088013725, `RNS_PRIME_BITS'd13242554, `RNS_PRIME_BITS'd1484483586, `RNS_PRIME_BITS'd687747905, `RNS_PRIME_BITS'd1165347914, `RNS_PRIME_BITS'd850830989, `RNS_PRIME_BITS'd179882299, `RNS_PRIME_BITS'd1100900306, `RNS_PRIME_BITS'd1898040454},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd965887127, `RNS_PRIME_BITS'd638065054, `RNS_PRIME_BITS'd944658461, `RNS_PRIME_BITS'd1003694775, `RNS_PRIME_BITS'd1348072526, `RNS_PRIME_BITS'd1888986692, `RNS_PRIME_BITS'd1248111520, `RNS_PRIME_BITS'd1318643875, `RNS_PRIME_BITS'd2137399927, `RNS_PRIME_BITS'd1483356111},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd901863058, `RNS_PRIME_BITS'd1697396893, `RNS_PRIME_BITS'd1332780340, `RNS_PRIME_BITS'd1033906560, `RNS_PRIME_BITS'd94672742, `RNS_PRIME_BITS'd1820774697, `RNS_PRIME_BITS'd1971389480, `RNS_PRIME_BITS'd1601738053, `RNS_PRIME_BITS'd669385788, `RNS_PRIME_BITS'd2078016371},
			'{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd708369181, `RNS_PRIME_BITS'd855258167, `RNS_PRIME_BITS'd208554435, `RNS_PRIME_BITS'd432078863, `RNS_PRIME_BITS'd1619495573, `RNS_PRIME_BITS'd1566689718, `RNS_PRIME_BITS'd813177745, `RNS_PRIME_BITS'd1315212570, `RNS_PRIME_BITS'd1421371015, `RNS_PRIME_BITS'd1175302112},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd2032375384, `RNS_PRIME_BITS'd153869869, `RNS_PRIME_BITS'd1114390586, `RNS_PRIME_BITS'd227929253, `RNS_PRIME_BITS'd1046230925, `RNS_PRIME_BITS'd960500751, `RNS_PRIME_BITS'd439426594, `RNS_PRIME_BITS'd1432117541, `RNS_PRIME_BITS'd647028451, `RNS_PRIME_BITS'd43125503},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd686368173, `RNS_PRIME_BITS'd1101027483, `RNS_PRIME_BITS'd1439990192, `RNS_PRIME_BITS'd1567734325, `RNS_PRIME_BITS'd1928804617, `RNS_PRIME_BITS'd759122739, `RNS_PRIME_BITS'd1664862721, `RNS_PRIME_BITS'd958354599, `RNS_PRIME_BITS'd628439079, `RNS_PRIME_BITS'd265280085},
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd1930745346, `RNS_PRIME_BITS'd1242643196, `RNS_PRIME_BITS'd931960151, `RNS_PRIME_BITS'd806838113, `RNS_PRIME_BITS'd1448017564, `RNS_PRIME_BITS'd1889291990, `RNS_PRIME_BITS'd174890120, `RNS_PRIME_BITS'd1405606306, `RNS_PRIME_BITS'd17299010, `RNS_PRIME_BITS'd1110613798},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd1223948152, `RNS_PRIME_BITS'd59750365, `RNS_PRIME_BITS'd824201308, `RNS_PRIME_BITS'd559292382, `RNS_PRIME_BITS'd1760010757, `RNS_PRIME_BITS'd715942105, `RNS_PRIME_BITS'd1731446105, `RNS_PRIME_BITS'd2131059015, `RNS_PRIME_BITS'd1923712156, `RNS_PRIME_BITS'd121855958},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd1422757924, `RNS_PRIME_BITS'd926677354, `RNS_PRIME_BITS'd1855196385, `RNS_PRIME_BITS'd1835021687, `RNS_PRIME_BITS'd1661608486, `RNS_PRIME_BITS'd1926377300, `RNS_PRIME_BITS'd651625814, `RNS_PRIME_BITS'd302993748, `RNS_PRIME_BITS'd1773741952, `RNS_PRIME_BITS'd1758363675},
			'{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd1832187758, `RNS_PRIME_BITS'd355263440, `RNS_PRIME_BITS'd230972645, `RNS_PRIME_BITS'd130058271, `RNS_PRIME_BITS'd1310586544, `RNS_PRIME_BITS'd20766307, `RNS_PRIME_BITS'd1608592228, `RNS_PRIME_BITS'd1267424663, `RNS_PRIME_BITS'd836425403, `RNS_PRIME_BITS'd165879156},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1512354342, `RNS_PRIME_BITS'd1214973053, `RNS_PRIME_BITS'd1134867455, `RNS_PRIME_BITS'd448105709, `RNS_PRIME_BITS'd1636078270, `RNS_PRIME_BITS'd1958061621, `RNS_PRIME_BITS'd2086671044, `RNS_PRIME_BITS'd1585104576, `RNS_PRIME_BITS'd1190630817, `RNS_PRIME_BITS'd1967138650},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd1966824096, `RNS_PRIME_BITS'd743527863, `RNS_PRIME_BITS'd1871248145, `RNS_PRIME_BITS'd1920799408, `RNS_PRIME_BITS'd1384075965, `RNS_PRIME_BITS'd1168359287, `RNS_PRIME_BITS'd1069821542, `RNS_PRIME_BITS'd1725878233, `RNS_PRIME_BITS'd157333049, `RNS_PRIME_BITS'd110870688},
			'{`RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd293939047, `RNS_PRIME_BITS'd89416979, `RNS_PRIME_BITS'd1711899231, `RNS_PRIME_BITS'd918333641, `RNS_PRIME_BITS'd699208034, `RNS_PRIME_BITS'd1337465825, `RNS_PRIME_BITS'd1176644344, `RNS_PRIME_BITS'd43454841, `RNS_PRIME_BITS'd1463992831, `RNS_PRIME_BITS'd1597042134},
			'{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd1358295062, `RNS_PRIME_BITS'd455625016, `RNS_PRIME_BITS'd866145584, `RNS_PRIME_BITS'd1037925824, `RNS_PRIME_BITS'd1436655550, `RNS_PRIME_BITS'd1195518986, `RNS_PRIME_BITS'd1610222772, `RNS_PRIME_BITS'd1817735815, `RNS_PRIME_BITS'd1269357152, `RNS_PRIME_BITS'd973317723},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd1224761672, `RNS_PRIME_BITS'd392345240, `RNS_PRIME_BITS'd1974190694, `RNS_PRIME_BITS'd1419316548, `RNS_PRIME_BITS'd753151536, `RNS_PRIME_BITS'd168287707, `RNS_PRIME_BITS'd602072643, `RNS_PRIME_BITS'd1417376311, `RNS_PRIME_BITS'd1148382389, `RNS_PRIME_BITS'd1732546477},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd1218272284, `RNS_PRIME_BITS'd1004833609, `RNS_PRIME_BITS'd1044859041, `RNS_PRIME_BITS'd873608925, `RNS_PRIME_BITS'd1186715704, `RNS_PRIME_BITS'd502189406, `RNS_PRIME_BITS'd2051404549, `RNS_PRIME_BITS'd239146010, `RNS_PRIME_BITS'd916771782, `RNS_PRIME_BITS'd1721612346},
			'{`RNS_PRIME_BITS'd132, `RNS_PRIME_BITS'd94966078, `RNS_PRIME_BITS'd1950500829, `RNS_PRIME_BITS'd312319856, `RNS_PRIME_BITS'd316226817, `RNS_PRIME_BITS'd1017312509, `RNS_PRIME_BITS'd513496360, `RNS_PRIME_BITS'd511752008, `RNS_PRIME_BITS'd960543387, `RNS_PRIME_BITS'd1876881962, `RNS_PRIME_BITS'd250426949},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd382366175, `RNS_PRIME_BITS'd840028000, `RNS_PRIME_BITS'd1380107556, `RNS_PRIME_BITS'd133957438, `RNS_PRIME_BITS'd1073552645, `RNS_PRIME_BITS'd1353475950, `RNS_PRIME_BITS'd1796365018, `RNS_PRIME_BITS'd470203826, `RNS_PRIME_BITS'd1699224200, `RNS_PRIME_BITS'd802388360},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd224509868, `RNS_PRIME_BITS'd1369742608, `RNS_PRIME_BITS'd455939089, `RNS_PRIME_BITS'd1032467332, `RNS_PRIME_BITS'd200974272, `RNS_PRIME_BITS'd604163912, `RNS_PRIME_BITS'd1649928229, `RNS_PRIME_BITS'd1546681827, `RNS_PRIME_BITS'd1156880120, `RNS_PRIME_BITS'd481966423},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd1818809183, `RNS_PRIME_BITS'd436311344, `RNS_PRIME_BITS'd272034618, `RNS_PRIME_BITS'd173580041, `RNS_PRIME_BITS'd1933231670, `RNS_PRIME_BITS'd1112203252, `RNS_PRIME_BITS'd1095445335, `RNS_PRIME_BITS'd744819199, `RNS_PRIME_BITS'd816531094, `RNS_PRIME_BITS'd1488434879},
			'{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd1727284613, `RNS_PRIME_BITS'd1806459492, `RNS_PRIME_BITS'd751494224, `RNS_PRIME_BITS'd1908934952, `RNS_PRIME_BITS'd1206892455, `RNS_PRIME_BITS'd1805501227, `RNS_PRIME_BITS'd424043786, `RNS_PRIME_BITS'd2045911239, `RNS_PRIME_BITS'd39062901, `RNS_PRIME_BITS'd2017185272},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1780981311, `RNS_PRIME_BITS'd809907616, `RNS_PRIME_BITS'd1442001684, `RNS_PRIME_BITS'd2039729648, `RNS_PRIME_BITS'd840657404, `RNS_PRIME_BITS'd1010149592, `RNS_PRIME_BITS'd1692689927, `RNS_PRIME_BITS'd1284498972, `RNS_PRIME_BITS'd141413674, `RNS_PRIME_BITS'd496895392},
			'{`RNS_PRIME_BITS'd66, `RNS_PRIME_BITS'd1460867205, `RNS_PRIME_BITS'd1963491127, `RNS_PRIME_BITS'd917452296, `RNS_PRIME_BITS'd1397652244, `RNS_PRIME_BITS'd1234474140, `RNS_PRIME_BITS'd1596901958, `RNS_PRIME_BITS'd1630203713, `RNS_PRIME_BITS'd1449924698, `RNS_PRIME_BITS'd1050091104, `RNS_PRIME_BITS'd820448346},
			'{`RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd1847241786, `RNS_PRIME_BITS'd341120682, `RNS_PRIME_BITS'd1652287903, `RNS_PRIME_BITS'd819352319, `RNS_PRIME_BITS'd1513853215, `RNS_PRIME_BITS'd1021877413, `RNS_PRIME_BITS'd1109033810, `RNS_PRIME_BITS'd1604018535, `RNS_PRIME_BITS'd1939458288, `RNS_PRIME_BITS'd1074272909},
			'{`RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd647789996, `RNS_PRIME_BITS'd573264143, `RNS_PRIME_BITS'd1902906456, `RNS_PRIME_BITS'd765882119, `RNS_PRIME_BITS'd1225986634, `RNS_PRIME_BITS'd1473111296, `RNS_PRIME_BITS'd707966785, `RNS_PRIME_BITS'd1043109791, `RNS_PRIME_BITS'd1358262689, `RNS_PRIME_BITS'd463388865}
		},
		'{
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd1830594593, `RNS_PRIME_BITS'd635052174, `RNS_PRIME_BITS'd1283010518, `RNS_PRIME_BITS'd1868454953, `RNS_PRIME_BITS'd1801455073, `RNS_PRIME_BITS'd308166474, `RNS_PRIME_BITS'd1517320037, `RNS_PRIME_BITS'd1448544719, `RNS_PRIME_BITS'd1929259717, `RNS_PRIME_BITS'd1751270350},
			'{`RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd471448206, `RNS_PRIME_BITS'd10284598, `RNS_PRIME_BITS'd2041542947, `RNS_PRIME_BITS'd1238665677, `RNS_PRIME_BITS'd912391353, `RNS_PRIME_BITS'd109072677, `RNS_PRIME_BITS'd1848597791, `RNS_PRIME_BITS'd132518041, `RNS_PRIME_BITS'd1097254034, `RNS_PRIME_BITS'd921031310},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd1595397622, `RNS_PRIME_BITS'd525003652, `RNS_PRIME_BITS'd1344430257, `RNS_PRIME_BITS'd1707330580, `RNS_PRIME_BITS'd300379262, `RNS_PRIME_BITS'd129079534, `RNS_PRIME_BITS'd812204283, `RNS_PRIME_BITS'd2311055, `RNS_PRIME_BITS'd227033748, `RNS_PRIME_BITS'd1915295557},
			'{`RNS_PRIME_BITS'd251, `RNS_PRIME_BITS'd1708907118, `RNS_PRIME_BITS'd617641436, `RNS_PRIME_BITS'd249632339, `RNS_PRIME_BITS'd818033043, `RNS_PRIME_BITS'd1479257858, `RNS_PRIME_BITS'd587042300, `RNS_PRIME_BITS'd458522204, `RNS_PRIME_BITS'd360485226, `RNS_PRIME_BITS'd2023623594, `RNS_PRIME_BITS'd775793888},
			'{`RNS_PRIME_BITS'd131, `RNS_PRIME_BITS'd769230889, `RNS_PRIME_BITS'd1946214386, `RNS_PRIME_BITS'd1657636874, `RNS_PRIME_BITS'd1444516340, `RNS_PRIME_BITS'd1833738462, `RNS_PRIME_BITS'd214620846, `RNS_PRIME_BITS'd1386822992, `RNS_PRIME_BITS'd41598877, `RNS_PRIME_BITS'd794730649, `RNS_PRIME_BITS'd1531723601},
			'{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd1597797665, `RNS_PRIME_BITS'd1146105962, `RNS_PRIME_BITS'd1663049317, `RNS_PRIME_BITS'd2074414179, `RNS_PRIME_BITS'd1603646855, `RNS_PRIME_BITS'd1452563860, `RNS_PRIME_BITS'd349271969, `RNS_PRIME_BITS'd1469279945, `RNS_PRIME_BITS'd891013558, `RNS_PRIME_BITS'd383308818},
			'{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd1092797308, `RNS_PRIME_BITS'd1308040833, `RNS_PRIME_BITS'd951601468, `RNS_PRIME_BITS'd1292775404, `RNS_PRIME_BITS'd2139045535, `RNS_PRIME_BITS'd1587067432, `RNS_PRIME_BITS'd38419700, `RNS_PRIME_BITS'd2097368885, `RNS_PRIME_BITS'd1546796792, `RNS_PRIME_BITS'd91558367},
			'{`RNS_PRIME_BITS'd244, `RNS_PRIME_BITS'd722168243, `RNS_PRIME_BITS'd1858757158, `RNS_PRIME_BITS'd543255036, `RNS_PRIME_BITS'd858285724, `RNS_PRIME_BITS'd813336374, `RNS_PRIME_BITS'd752218571, `RNS_PRIME_BITS'd180607074, `RNS_PRIME_BITS'd1267038139, `RNS_PRIME_BITS'd600719418, `RNS_PRIME_BITS'd286088174},
			'{`RNS_PRIME_BITS'd140, `RNS_PRIME_BITS'd1099102855, `RNS_PRIME_BITS'd275496277, `RNS_PRIME_BITS'd107900356, `RNS_PRIME_BITS'd1192759325, `RNS_PRIME_BITS'd987618330, `RNS_PRIME_BITS'd934761993, `RNS_PRIME_BITS'd1156696837, `RNS_PRIME_BITS'd1869619114, `RNS_PRIME_BITS'd1607159737, `RNS_PRIME_BITS'd1025719108},
			'{`RNS_PRIME_BITS'd209, `RNS_PRIME_BITS'd63464056, `RNS_PRIME_BITS'd1750884091, `RNS_PRIME_BITS'd1329595715, `RNS_PRIME_BITS'd1940196449, `RNS_PRIME_BITS'd1972400413, `RNS_PRIME_BITS'd1757726183, `RNS_PRIME_BITS'd276839822, `RNS_PRIME_BITS'd1037223245, `RNS_PRIME_BITS'd2118865000, `RNS_PRIME_BITS'd272451573},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd75082068, `RNS_PRIME_BITS'd1387989277, `RNS_PRIME_BITS'd1755308462, `RNS_PRIME_BITS'd1216142778, `RNS_PRIME_BITS'd1352705718, `RNS_PRIME_BITS'd258022345, `RNS_PRIME_BITS'd1331050810, `RNS_PRIME_BITS'd1581778185, `RNS_PRIME_BITS'd1473036566, `RNS_PRIME_BITS'd1647433610},
			'{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd1864192010, `RNS_PRIME_BITS'd1016777977, `RNS_PRIME_BITS'd1921798665, `RNS_PRIME_BITS'd1872859260, `RNS_PRIME_BITS'd1067932573, `RNS_PRIME_BITS'd1558761174, `RNS_PRIME_BITS'd1557375120, `RNS_PRIME_BITS'd1183222752, `RNS_PRIME_BITS'd1125554427, `RNS_PRIME_BITS'd1246882625},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd1754398022, `RNS_PRIME_BITS'd1989463697, `RNS_PRIME_BITS'd1395292099, `RNS_PRIME_BITS'd1204873373, `RNS_PRIME_BITS'd139681625, `RNS_PRIME_BITS'd654497065, `RNS_PRIME_BITS'd2039430311, `RNS_PRIME_BITS'd635754057, `RNS_PRIME_BITS'd509727324, `RNS_PRIME_BITS'd1896536073},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd839238125, `RNS_PRIME_BITS'd1469507393, `RNS_PRIME_BITS'd1782531712, `RNS_PRIME_BITS'd909549490, `RNS_PRIME_BITS'd382941012, `RNS_PRIME_BITS'd1876973435, `RNS_PRIME_BITS'd1620381764, `RNS_PRIME_BITS'd1605205471, `RNS_PRIME_BITS'd136321693, `RNS_PRIME_BITS'd1549535846},
			'{`RNS_PRIME_BITS'd148, `RNS_PRIME_BITS'd1354528461, `RNS_PRIME_BITS'd1611051046, `RNS_PRIME_BITS'd199071660, `RNS_PRIME_BITS'd437110477, `RNS_PRIME_BITS'd1157127670, `RNS_PRIME_BITS'd2039532777, `RNS_PRIME_BITS'd545963928, `RNS_PRIME_BITS'd1127376740, `RNS_PRIME_BITS'd1376003511, `RNS_PRIME_BITS'd1745933575},
			'{`RNS_PRIME_BITS'd147, `RNS_PRIME_BITS'd54307582, `RNS_PRIME_BITS'd294106283, `RNS_PRIME_BITS'd1222799633, `RNS_PRIME_BITS'd895184227, `RNS_PRIME_BITS'd494448735, `RNS_PRIME_BITS'd589602968, `RNS_PRIME_BITS'd273122676, `RNS_PRIME_BITS'd1340090172, `RNS_PRIME_BITS'd151827560, `RNS_PRIME_BITS'd1814996861},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd1830900760, `RNS_PRIME_BITS'd793234455, `RNS_PRIME_BITS'd1480319799, `RNS_PRIME_BITS'd1428979957, `RNS_PRIME_BITS'd716220952, `RNS_PRIME_BITS'd440348454, `RNS_PRIME_BITS'd1550485207, `RNS_PRIME_BITS'd1117715500, `RNS_PRIME_BITS'd620964777, `RNS_PRIME_BITS'd614983979},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd45474555, `RNS_PRIME_BITS'd200160850, `RNS_PRIME_BITS'd875308062, `RNS_PRIME_BITS'd1456739501, `RNS_PRIME_BITS'd1289441699, `RNS_PRIME_BITS'd2083488080, `RNS_PRIME_BITS'd1990230137, `RNS_PRIME_BITS'd1247146457, `RNS_PRIME_BITS'd1203120989, `RNS_PRIME_BITS'd821376191},
			'{`RNS_PRIME_BITS'd179, `RNS_PRIME_BITS'd2009040287, `RNS_PRIME_BITS'd2119258449, `RNS_PRIME_BITS'd705780947, `RNS_PRIME_BITS'd1305566096, `RNS_PRIME_BITS'd368642947, `RNS_PRIME_BITS'd1766833568, `RNS_PRIME_BITS'd323069027, `RNS_PRIME_BITS'd1611977621, `RNS_PRIME_BITS'd625170064, `RNS_PRIME_BITS'd209191650},
			'{`RNS_PRIME_BITS'd254, `RNS_PRIME_BITS'd27324387, `RNS_PRIME_BITS'd80862483, `RNS_PRIME_BITS'd1107881401, `RNS_PRIME_BITS'd1893344701, `RNS_PRIME_BITS'd1298058012, `RNS_PRIME_BITS'd650407461, `RNS_PRIME_BITS'd165965186, `RNS_PRIME_BITS'd161513798, `RNS_PRIME_BITS'd983088889, `RNS_PRIME_BITS'd318460599},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd1149540269, `RNS_PRIME_BITS'd1303347717, `RNS_PRIME_BITS'd674815698, `RNS_PRIME_BITS'd840619572, `RNS_PRIME_BITS'd92175099, `RNS_PRIME_BITS'd1065373451, `RNS_PRIME_BITS'd366624196, `RNS_PRIME_BITS'd1799646045, `RNS_PRIME_BITS'd1123767382, `RNS_PRIME_BITS'd1662999417},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd1722519682, `RNS_PRIME_BITS'd1314612176, `RNS_PRIME_BITS'd1819646102, `RNS_PRIME_BITS'd482409380, `RNS_PRIME_BITS'd1887509616, `RNS_PRIME_BITS'd344164170, `RNS_PRIME_BITS'd1854183272, `RNS_PRIME_BITS'd1899904035, `RNS_PRIME_BITS'd785414278, `RNS_PRIME_BITS'd196751530},
			'{`RNS_PRIME_BITS'd179, `RNS_PRIME_BITS'd1171284569, `RNS_PRIME_BITS'd1739118080, `RNS_PRIME_BITS'd225129441, `RNS_PRIME_BITS'd1779589231, `RNS_PRIME_BITS'd9363896, `RNS_PRIME_BITS'd1624126486, `RNS_PRIME_BITS'd2116796999, `RNS_PRIME_BITS'd1264463887, `RNS_PRIME_BITS'd1181322318, `RNS_PRIME_BITS'd589964074},
			'{`RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd1480362259, `RNS_PRIME_BITS'd1336311897, `RNS_PRIME_BITS'd849305081, `RNS_PRIME_BITS'd689246040, `RNS_PRIME_BITS'd686454469, `RNS_PRIME_BITS'd1237071807, `RNS_PRIME_BITS'd930555815, `RNS_PRIME_BITS'd473627697, `RNS_PRIME_BITS'd1866113568, `RNS_PRIME_BITS'd853570649},
			'{`RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd1430356764, `RNS_PRIME_BITS'd855269182, `RNS_PRIME_BITS'd1355923164, `RNS_PRIME_BITS'd1515380931, `RNS_PRIME_BITS'd356622209, `RNS_PRIME_BITS'd2075467109, `RNS_PRIME_BITS'd297352735, `RNS_PRIME_BITS'd590617367, `RNS_PRIME_BITS'd309638650, `RNS_PRIME_BITS'd1196795586},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1283284787, `RNS_PRIME_BITS'd726548834, `RNS_PRIME_BITS'd1701790351, `RNS_PRIME_BITS'd665740836, `RNS_PRIME_BITS'd184774413, `RNS_PRIME_BITS'd912046426, `RNS_PRIME_BITS'd4229079, `RNS_PRIME_BITS'd1320229163, `RNS_PRIME_BITS'd1097524966, `RNS_PRIME_BITS'd983256081},
			'{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd203015582, `RNS_PRIME_BITS'd143165313, `RNS_PRIME_BITS'd466498958, `RNS_PRIME_BITS'd1001447576, `RNS_PRIME_BITS'd1618424708, `RNS_PRIME_BITS'd424232457, `RNS_PRIME_BITS'd817152424, `RNS_PRIME_BITS'd1250457628, `RNS_PRIME_BITS'd594249455, `RNS_PRIME_BITS'd529138325},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd1375235903, `RNS_PRIME_BITS'd683237374, `RNS_PRIME_BITS'd1342170533, `RNS_PRIME_BITS'd2134842792, `RNS_PRIME_BITS'd1272653185, `RNS_PRIME_BITS'd662734736, `RNS_PRIME_BITS'd331417844, `RNS_PRIME_BITS'd1249548740, `RNS_PRIME_BITS'd1558779015, `RNS_PRIME_BITS'd1862418350},
			'{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd227461782, `RNS_PRIME_BITS'd1192047266, `RNS_PRIME_BITS'd1436040955, `RNS_PRIME_BITS'd1960525897, `RNS_PRIME_BITS'd1474722258, `RNS_PRIME_BITS'd1235373487, `RNS_PRIME_BITS'd1353648216, `RNS_PRIME_BITS'd590614606, `RNS_PRIME_BITS'd288809502, `RNS_PRIME_BITS'd546751118},
			'{`RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd1150362782, `RNS_PRIME_BITS'd368606169, `RNS_PRIME_BITS'd1859167521, `RNS_PRIME_BITS'd584616639, `RNS_PRIME_BITS'd2059284756, `RNS_PRIME_BITS'd55990657, `RNS_PRIME_BITS'd2035917418, `RNS_PRIME_BITS'd1439322006, `RNS_PRIME_BITS'd1048846475, `RNS_PRIME_BITS'd707904313},
			'{`RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd1931095045, `RNS_PRIME_BITS'd1476319930, `RNS_PRIME_BITS'd1086597405, `RNS_PRIME_BITS'd1702908355, `RNS_PRIME_BITS'd493403952, `RNS_PRIME_BITS'd625879920, `RNS_PRIME_BITS'd704910542, `RNS_PRIME_BITS'd233630602, `RNS_PRIME_BITS'd1605274830, `RNS_PRIME_BITS'd95154695},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1239255884, `RNS_PRIME_BITS'd1617373145, `RNS_PRIME_BITS'd1791972888, `RNS_PRIME_BITS'd1135359336, `RNS_PRIME_BITS'd1915162756, `RNS_PRIME_BITS'd1468542201, `RNS_PRIME_BITS'd1031551067, `RNS_PRIME_BITS'd59976946, `RNS_PRIME_BITS'd1299333287, `RNS_PRIME_BITS'd1540488650},
			'{`RNS_PRIME_BITS'd108, `RNS_PRIME_BITS'd152104724, `RNS_PRIME_BITS'd1469823516, `RNS_PRIME_BITS'd698173873, `RNS_PRIME_BITS'd1410165174, `RNS_PRIME_BITS'd604889259, `RNS_PRIME_BITS'd1540847599, `RNS_PRIME_BITS'd2014187173, `RNS_PRIME_BITS'd425715105, `RNS_PRIME_BITS'd1772138011, `RNS_PRIME_BITS'd151182488},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd2073690772, `RNS_PRIME_BITS'd1980839883, `RNS_PRIME_BITS'd1164381351, `RNS_PRIME_BITS'd1505981619, `RNS_PRIME_BITS'd979036372, `RNS_PRIME_BITS'd586147271, `RNS_PRIME_BITS'd1597829504, `RNS_PRIME_BITS'd1275517068, `RNS_PRIME_BITS'd1282592903, `RNS_PRIME_BITS'd985192939},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd1083086377, `RNS_PRIME_BITS'd1885322725, `RNS_PRIME_BITS'd1227246667, `RNS_PRIME_BITS'd164558840, `RNS_PRIME_BITS'd785846137, `RNS_PRIME_BITS'd1638964343, `RNS_PRIME_BITS'd353148682, `RNS_PRIME_BITS'd1739493258, `RNS_PRIME_BITS'd957636840, `RNS_PRIME_BITS'd338139443},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd236115242, `RNS_PRIME_BITS'd1605658973, `RNS_PRIME_BITS'd1089256958, `RNS_PRIME_BITS'd260461459, `RNS_PRIME_BITS'd668884049, `RNS_PRIME_BITS'd430366057, `RNS_PRIME_BITS'd843943309, `RNS_PRIME_BITS'd408124808, `RNS_PRIME_BITS'd1957739356, `RNS_PRIME_BITS'd165973560},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd816046015, `RNS_PRIME_BITS'd358020963, `RNS_PRIME_BITS'd1209107465, `RNS_PRIME_BITS'd1159748344, `RNS_PRIME_BITS'd2045427214, `RNS_PRIME_BITS'd170582553, `RNS_PRIME_BITS'd323938533, `RNS_PRIME_BITS'd408680801, `RNS_PRIME_BITS'd1128417752, `RNS_PRIME_BITS'd896880240},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1817067578, `RNS_PRIME_BITS'd1894790006, `RNS_PRIME_BITS'd2001175412, `RNS_PRIME_BITS'd425659546, `RNS_PRIME_BITS'd2052025236, `RNS_PRIME_BITS'd1855095080, `RNS_PRIME_BITS'd1364871431, `RNS_PRIME_BITS'd995571920, `RNS_PRIME_BITS'd1334870089, `RNS_PRIME_BITS'd1955567284},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1815993801, `RNS_PRIME_BITS'd295921616, `RNS_PRIME_BITS'd1192258502, `RNS_PRIME_BITS'd714583703, `RNS_PRIME_BITS'd267919233, `RNS_PRIME_BITS'd594209386, `RNS_PRIME_BITS'd1923614236, `RNS_PRIME_BITS'd574613333, `RNS_PRIME_BITS'd1809368510, `RNS_PRIME_BITS'd776646878},
			'{`RNS_PRIME_BITS'd250, `RNS_PRIME_BITS'd203319519, `RNS_PRIME_BITS'd523307638, `RNS_PRIME_BITS'd1446234699, `RNS_PRIME_BITS'd2118127220, `RNS_PRIME_BITS'd1649919456, `RNS_PRIME_BITS'd1370963151, `RNS_PRIME_BITS'd1367672864, `RNS_PRIME_BITS'd78818034, `RNS_PRIME_BITS'd1901131716, `RNS_PRIME_BITS'd848377944},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd322291579, `RNS_PRIME_BITS'd1895029670, `RNS_PRIME_BITS'd1683638941, `RNS_PRIME_BITS'd1778212760, `RNS_PRIME_BITS'd1943895310, `RNS_PRIME_BITS'd1596476809, `RNS_PRIME_BITS'd1027715214, `RNS_PRIME_BITS'd1025088437, `RNS_PRIME_BITS'd1427850875, `RNS_PRIME_BITS'd797650963},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd835630192, `RNS_PRIME_BITS'd1514398200, `RNS_PRIME_BITS'd691644903, `RNS_PRIME_BITS'd1962727006, `RNS_PRIME_BITS'd422117785, `RNS_PRIME_BITS'd731891235, `RNS_PRIME_BITS'd1547850339, `RNS_PRIME_BITS'd1585518753, `RNS_PRIME_BITS'd246250761, `RNS_PRIME_BITS'd1559492797},
			'{`RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd2025360953, `RNS_PRIME_BITS'd97707405, `RNS_PRIME_BITS'd1407933586, `RNS_PRIME_BITS'd2097009987, `RNS_PRIME_BITS'd2060702414, `RNS_PRIME_BITS'd720016146, `RNS_PRIME_BITS'd414936042, `RNS_PRIME_BITS'd161641320, `RNS_PRIME_BITS'd1532729583, `RNS_PRIME_BITS'd1187273283},
			'{`RNS_PRIME_BITS'd154, `RNS_PRIME_BITS'd575630178, `RNS_PRIME_BITS'd782551085, `RNS_PRIME_BITS'd800307106, `RNS_PRIME_BITS'd360972388, `RNS_PRIME_BITS'd1865980170, `RNS_PRIME_BITS'd1768020781, `RNS_PRIME_BITS'd1154217848, `RNS_PRIME_BITS'd396856914, `RNS_PRIME_BITS'd126558609, `RNS_PRIME_BITS'd1106886637},
			'{`RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd938033732, `RNS_PRIME_BITS'd1418183847, `RNS_PRIME_BITS'd1836226493, `RNS_PRIME_BITS'd202581803, `RNS_PRIME_BITS'd827957282, `RNS_PRIME_BITS'd1320164473, `RNS_PRIME_BITS'd568452565, `RNS_PRIME_BITS'd1332781154, `RNS_PRIME_BITS'd972276663, `RNS_PRIME_BITS'd1764674617},
			'{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd1746679769, `RNS_PRIME_BITS'd226967150, `RNS_PRIME_BITS'd478593949, `RNS_PRIME_BITS'd1739154617, `RNS_PRIME_BITS'd33793707, `RNS_PRIME_BITS'd1929839264, `RNS_PRIME_BITS'd406738871, `RNS_PRIME_BITS'd247919767, `RNS_PRIME_BITS'd592619974, `RNS_PRIME_BITS'd1821460386},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd1273101156, `RNS_PRIME_BITS'd397569435, `RNS_PRIME_BITS'd420131109, `RNS_PRIME_BITS'd1381067359, `RNS_PRIME_BITS'd2045165831, `RNS_PRIME_BITS'd858666945, `RNS_PRIME_BITS'd238159785, `RNS_PRIME_BITS'd774328045, `RNS_PRIME_BITS'd1223675914, `RNS_PRIME_BITS'd1012568179},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd250619387, `RNS_PRIME_BITS'd1942540011, `RNS_PRIME_BITS'd1295784651, `RNS_PRIME_BITS'd2061731676, `RNS_PRIME_BITS'd1674296503, `RNS_PRIME_BITS'd174551035, `RNS_PRIME_BITS'd885281242, `RNS_PRIME_BITS'd620570659, `RNS_PRIME_BITS'd2112337508, `RNS_PRIME_BITS'd1705186646},
			'{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd1487391608, `RNS_PRIME_BITS'd1106953801, `RNS_PRIME_BITS'd920384915, `RNS_PRIME_BITS'd1062406747, `RNS_PRIME_BITS'd1083643074, `RNS_PRIME_BITS'd1260726341, `RNS_PRIME_BITS'd690944159, `RNS_PRIME_BITS'd384751918, `RNS_PRIME_BITS'd2026292886, `RNS_PRIME_BITS'd842984813},
			'{`RNS_PRIME_BITS'd33, `RNS_PRIME_BITS'd1933355743, `RNS_PRIME_BITS'd906508753, `RNS_PRIME_BITS'd1382142376, `RNS_PRIME_BITS'd1573273505, `RNS_PRIME_BITS'd828993086, `RNS_PRIME_BITS'd2069897245, `RNS_PRIME_BITS'd1107644755, `RNS_PRIME_BITS'd1847562376, `RNS_PRIME_BITS'd2136088163, `RNS_PRIME_BITS'd2089601301},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd1987405791, `RNS_PRIME_BITS'd751577849, `RNS_PRIME_BITS'd106817608, `RNS_PRIME_BITS'd1928338662, `RNS_PRIME_BITS'd609330356, `RNS_PRIME_BITS'd706564875, `RNS_PRIME_BITS'd852565921, `RNS_PRIME_BITS'd190150785, `RNS_PRIME_BITS'd1301586875, `RNS_PRIME_BITS'd1139528448},
			'{`RNS_PRIME_BITS'd167, `RNS_PRIME_BITS'd67500971, `RNS_PRIME_BITS'd1391130517, `RNS_PRIME_BITS'd484149956, `RNS_PRIME_BITS'd568707576, `RNS_PRIME_BITS'd867639538, `RNS_PRIME_BITS'd1909766520, `RNS_PRIME_BITS'd1621328526, `RNS_PRIME_BITS'd858338612, `RNS_PRIME_BITS'd285596872, `RNS_PRIME_BITS'd210455881},
			'{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd1850565286, `RNS_PRIME_BITS'd2027159529, `RNS_PRIME_BITS'd279761875, `RNS_PRIME_BITS'd786677892, `RNS_PRIME_BITS'd1707795165, `RNS_PRIME_BITS'd1516542895, `RNS_PRIME_BITS'd1826162517, `RNS_PRIME_BITS'd1793610089, `RNS_PRIME_BITS'd1559151262, `RNS_PRIME_BITS'd688343551},
			'{`RNS_PRIME_BITS'd180, `RNS_PRIME_BITS'd1105260684, `RNS_PRIME_BITS'd28546864, `RNS_PRIME_BITS'd1054790336, `RNS_PRIME_BITS'd1459218005, `RNS_PRIME_BITS'd845528046, `RNS_PRIME_BITS'd589782325, `RNS_PRIME_BITS'd1373769191, `RNS_PRIME_BITS'd1837367445, `RNS_PRIME_BITS'd136486927, `RNS_PRIME_BITS'd697541219},
			'{`RNS_PRIME_BITS'd108, `RNS_PRIME_BITS'd390630714, `RNS_PRIME_BITS'd950840355, `RNS_PRIME_BITS'd1856098391, `RNS_PRIME_BITS'd2091506787, `RNS_PRIME_BITS'd950676547, `RNS_PRIME_BITS'd1188169689, `RNS_PRIME_BITS'd2139975840, `RNS_PRIME_BITS'd1054929471, `RNS_PRIME_BITS'd1920281639, `RNS_PRIME_BITS'd761632005},
			'{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd825457133, `RNS_PRIME_BITS'd1580961986, `RNS_PRIME_BITS'd1522978897, `RNS_PRIME_BITS'd1986747765, `RNS_PRIME_BITS'd179456863, `RNS_PRIME_BITS'd1986888053, `RNS_PRIME_BITS'd303849609, `RNS_PRIME_BITS'd657232242, `RNS_PRIME_BITS'd1713743417, `RNS_PRIME_BITS'd842682303},
			'{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd1877260669, `RNS_PRIME_BITS'd600387412, `RNS_PRIME_BITS'd1849669741, `RNS_PRIME_BITS'd1589193400, `RNS_PRIME_BITS'd1651565532, `RNS_PRIME_BITS'd1335176854, `RNS_PRIME_BITS'd1036912402, `RNS_PRIME_BITS'd734694377, `RNS_PRIME_BITS'd879145868, `RNS_PRIME_BITS'd1563888499},
			'{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd2031517891, `RNS_PRIME_BITS'd1468023818, `RNS_PRIME_BITS'd2115606989, `RNS_PRIME_BITS'd834168729, `RNS_PRIME_BITS'd1498930860, `RNS_PRIME_BITS'd297110765, `RNS_PRIME_BITS'd2026451118, `RNS_PRIME_BITS'd1750783798, `RNS_PRIME_BITS'd1527701202, `RNS_PRIME_BITS'd2073460895},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd1204542843, `RNS_PRIME_BITS'd431209017, `RNS_PRIME_BITS'd1297460400, `RNS_PRIME_BITS'd304253696, `RNS_PRIME_BITS'd2113793015, `RNS_PRIME_BITS'd195051616, `RNS_PRIME_BITS'd1660027936, `RNS_PRIME_BITS'd1012701290, `RNS_PRIME_BITS'd1730437683, `RNS_PRIME_BITS'd603216054},
			'{`RNS_PRIME_BITS'd43, `RNS_PRIME_BITS'd1321157133, `RNS_PRIME_BITS'd1628537374, `RNS_PRIME_BITS'd529481590, `RNS_PRIME_BITS'd14123723, `RNS_PRIME_BITS'd1236211715, `RNS_PRIME_BITS'd288145560, `RNS_PRIME_BITS'd1368002439, `RNS_PRIME_BITS'd196365195, `RNS_PRIME_BITS'd1793059820, `RNS_PRIME_BITS'd171907509},
			'{`RNS_PRIME_BITS'd93, `RNS_PRIME_BITS'd1495439818, `RNS_PRIME_BITS'd1955014566, `RNS_PRIME_BITS'd51902079, `RNS_PRIME_BITS'd1271107478, `RNS_PRIME_BITS'd1522751221, `RNS_PRIME_BITS'd1669310722, `RNS_PRIME_BITS'd574123812, `RNS_PRIME_BITS'd771168349, `RNS_PRIME_BITS'd2136222284, `RNS_PRIME_BITS'd1782063075},
			'{`RNS_PRIME_BITS'd138, `RNS_PRIME_BITS'd102646347, `RNS_PRIME_BITS'd207023397, `RNS_PRIME_BITS'd1446956487, `RNS_PRIME_BITS'd692499020, `RNS_PRIME_BITS'd1302377048, `RNS_PRIME_BITS'd1051505232, `RNS_PRIME_BITS'd87973492, `RNS_PRIME_BITS'd1534564311, `RNS_PRIME_BITS'd1941235508, `RNS_PRIME_BITS'd1538251482},
			'{`RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd664852889, `RNS_PRIME_BITS'd1167490248, `RNS_PRIME_BITS'd552628490, `RNS_PRIME_BITS'd542136375, `RNS_PRIME_BITS'd947520481, `RNS_PRIME_BITS'd113833946, `RNS_PRIME_BITS'd1951856509, `RNS_PRIME_BITS'd1749185018, `RNS_PRIME_BITS'd685799117, `RNS_PRIME_BITS'd1813914150},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd1107186936, `RNS_PRIME_BITS'd1940302764, `RNS_PRIME_BITS'd1939581998, `RNS_PRIME_BITS'd951940249, `RNS_PRIME_BITS'd1369339996, `RNS_PRIME_BITS'd1263987944, `RNS_PRIME_BITS'd1131072564, `RNS_PRIME_BITS'd1798966457, `RNS_PRIME_BITS'd431790400, `RNS_PRIME_BITS'd657139696}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd1894736973, `RNS_PRIME_BITS'd784217465, `RNS_PRIME_BITS'd2038291888, `RNS_PRIME_BITS'd1716956691, `RNS_PRIME_BITS'd1752673844, `RNS_PRIME_BITS'd1854126027, `RNS_PRIME_BITS'd2098968497, `RNS_PRIME_BITS'd1741520124, `RNS_PRIME_BITS'd1789768460, `RNS_PRIME_BITS'd212309001},
			'{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd2031348663, `RNS_PRIME_BITS'd1927675409, `RNS_PRIME_BITS'd203376966, `RNS_PRIME_BITS'd1055582093, `RNS_PRIME_BITS'd1527705661, `RNS_PRIME_BITS'd1382356666, `RNS_PRIME_BITS'd1546242777, `RNS_PRIME_BITS'd728667211, `RNS_PRIME_BITS'd2019048699, `RNS_PRIME_BITS'd734017170},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd1398718732, `RNS_PRIME_BITS'd1803042816, `RNS_PRIME_BITS'd844265329, `RNS_PRIME_BITS'd81610673, `RNS_PRIME_BITS'd559307702, `RNS_PRIME_BITS'd355382446, `RNS_PRIME_BITS'd1354603284, `RNS_PRIME_BITS'd370239913, `RNS_PRIME_BITS'd934841153, `RNS_PRIME_BITS'd1897500022},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd2088885210, `RNS_PRIME_BITS'd1805162228, `RNS_PRIME_BITS'd2047394668, `RNS_PRIME_BITS'd1711459801, `RNS_PRIME_BITS'd1541158891, `RNS_PRIME_BITS'd2094120779, `RNS_PRIME_BITS'd117160621, `RNS_PRIME_BITS'd1493600233, `RNS_PRIME_BITS'd110502899, `RNS_PRIME_BITS'd656753225},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd1122998748, `RNS_PRIME_BITS'd625830662, `RNS_PRIME_BITS'd388113819, `RNS_PRIME_BITS'd2035390491, `RNS_PRIME_BITS'd713259247, `RNS_PRIME_BITS'd1194438850, `RNS_PRIME_BITS'd1964580646, `RNS_PRIME_BITS'd1530347451, `RNS_PRIME_BITS'd882221572, `RNS_PRIME_BITS'd2125503037},
			'{`RNS_PRIME_BITS'd63, `RNS_PRIME_BITS'd928017860, `RNS_PRIME_BITS'd142786996, `RNS_PRIME_BITS'd127046322, `RNS_PRIME_BITS'd808771334, `RNS_PRIME_BITS'd1676104489, `RNS_PRIME_BITS'd1572345723, `RNS_PRIME_BITS'd1438043398, `RNS_PRIME_BITS'd1069101662, `RNS_PRIME_BITS'd1958721293, `RNS_PRIME_BITS'd19726431},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd365687374, `RNS_PRIME_BITS'd1180186395, `RNS_PRIME_BITS'd855563579, `RNS_PRIME_BITS'd2002377631, `RNS_PRIME_BITS'd1987112191, `RNS_PRIME_BITS'd1003842129, `RNS_PRIME_BITS'd1741424702, `RNS_PRIME_BITS'd1620807945, `RNS_PRIME_BITS'd1870415188, `RNS_PRIME_BITS'd94338220},
			'{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd1481546344, `RNS_PRIME_BITS'd1750766142, `RNS_PRIME_BITS'd455267761, `RNS_PRIME_BITS'd1426011701, `RNS_PRIME_BITS'd2080412029, `RNS_PRIME_BITS'd790829049, `RNS_PRIME_BITS'd2067877069, `RNS_PRIME_BITS'd673787331, `RNS_PRIME_BITS'd1873357003, `RNS_PRIME_BITS'd1188025713},
			'{`RNS_PRIME_BITS'd252, `RNS_PRIME_BITS'd1574415978, `RNS_PRIME_BITS'd402877308, `RNS_PRIME_BITS'd872148956, `RNS_PRIME_BITS'd939014429, `RNS_PRIME_BITS'd1853902700, `RNS_PRIME_BITS'd1356356420, `RNS_PRIME_BITS'd343630257, `RNS_PRIME_BITS'd1723988937, `RNS_PRIME_BITS'd1631326364, `RNS_PRIME_BITS'd1693568215},
			'{`RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd1828329262, `RNS_PRIME_BITS'd1231613327, `RNS_PRIME_BITS'd1794974621, `RNS_PRIME_BITS'd1510801179, `RNS_PRIME_BITS'd428364426, `RNS_PRIME_BITS'd1178120200, `RNS_PRIME_BITS'd1364286401, `RNS_PRIME_BITS'd1550539376, `RNS_PRIME_BITS'd1264270463, `RNS_PRIME_BITS'd329042924},
			'{`RNS_PRIME_BITS'd109, `RNS_PRIME_BITS'd1721767427, `RNS_PRIME_BITS'd719080628, `RNS_PRIME_BITS'd349864445, `RNS_PRIME_BITS'd1164274416, `RNS_PRIME_BITS'd915072584, `RNS_PRIME_BITS'd944008541, `RNS_PRIME_BITS'd522854153, `RNS_PRIME_BITS'd1600478588, `RNS_PRIME_BITS'd2056363618, `RNS_PRIME_BITS'd897601035},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd2079582940, `RNS_PRIME_BITS'd1525173856, `RNS_PRIME_BITS'd1292243466, `RNS_PRIME_BITS'd1911587549, `RNS_PRIME_BITS'd1094505838, `RNS_PRIME_BITS'd1174963477, `RNS_PRIME_BITS'd829342937, `RNS_PRIME_BITS'd188252983, `RNS_PRIME_BITS'd1022324081, `RNS_PRIME_BITS'd1018314988},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd2011568867, `RNS_PRIME_BITS'd767794497, `RNS_PRIME_BITS'd2135051953, `RNS_PRIME_BITS'd1370615671, `RNS_PRIME_BITS'd179337303, `RNS_PRIME_BITS'd1357952016, `RNS_PRIME_BITS'd618482488, `RNS_PRIME_BITS'd639339809, `RNS_PRIME_BITS'd1273888863, `RNS_PRIME_BITS'd1997108103},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd1319020715, `RNS_PRIME_BITS'd603907508, `RNS_PRIME_BITS'd2013786546, `RNS_PRIME_BITS'd260768423, `RNS_PRIME_BITS'd1535838563, `RNS_PRIME_BITS'd1545958402, `RNS_PRIME_BITS'd168254335, `RNS_PRIME_BITS'd870357026, `RNS_PRIME_BITS'd1848337960, `RNS_PRIME_BITS'd579301844},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd762833733, `RNS_PRIME_BITS'd1616034882, `RNS_PRIME_BITS'd774937267, `RNS_PRIME_BITS'd1101600704, `RNS_PRIME_BITS'd840917968, `RNS_PRIME_BITS'd840626784, `RNS_PRIME_BITS'd1406269015, `RNS_PRIME_BITS'd688849970, `RNS_PRIME_BITS'd1001240806, `RNS_PRIME_BITS'd907528979},
			'{`RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd1985917159, `RNS_PRIME_BITS'd1266721215, `RNS_PRIME_BITS'd485383343, `RNS_PRIME_BITS'd805162661, `RNS_PRIME_BITS'd1383325834, `RNS_PRIME_BITS'd2067160420, `RNS_PRIME_BITS'd956652373, `RNS_PRIME_BITS'd1225748689, `RNS_PRIME_BITS'd871244966, `RNS_PRIME_BITS'd1048543595},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd1055040398, `RNS_PRIME_BITS'd978303215, `RNS_PRIME_BITS'd1256981549, `RNS_PRIME_BITS'd1904176916, `RNS_PRIME_BITS'd891503333, `RNS_PRIME_BITS'd1749763825, `RNS_PRIME_BITS'd668628743, `RNS_PRIME_BITS'd2074558391, `RNS_PRIME_BITS'd19828557, `RNS_PRIME_BITS'd1054139503},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd579179537, `RNS_PRIME_BITS'd866234750, `RNS_PRIME_BITS'd651979073, `RNS_PRIME_BITS'd835782282, `RNS_PRIME_BITS'd455963313, `RNS_PRIME_BITS'd1046023719, `RNS_PRIME_BITS'd82811289, `RNS_PRIME_BITS'd1662126254, `RNS_PRIME_BITS'd404110894, `RNS_PRIME_BITS'd1324495362},
			'{`RNS_PRIME_BITS'd12, `RNS_PRIME_BITS'd1394574200, `RNS_PRIME_BITS'd1529629882, `RNS_PRIME_BITS'd722907224, `RNS_PRIME_BITS'd957169463, `RNS_PRIME_BITS'd65489569, `RNS_PRIME_BITS'd2012361196, `RNS_PRIME_BITS'd1857940664, `RNS_PRIME_BITS'd1721452603, `RNS_PRIME_BITS'd967561577, `RNS_PRIME_BITS'd1332803573},
			'{`RNS_PRIME_BITS'd125, `RNS_PRIME_BITS'd602071633, `RNS_PRIME_BITS'd442739792, `RNS_PRIME_BITS'd77740530, `RNS_PRIME_BITS'd1839550137, `RNS_PRIME_BITS'd1613482433, `RNS_PRIME_BITS'd285728457, `RNS_PRIME_BITS'd898592314, `RNS_PRIME_BITS'd1021653282, `RNS_PRIME_BITS'd1751753272, `RNS_PRIME_BITS'd1539419869},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd851928034, `RNS_PRIME_BITS'd1515898945, `RNS_PRIME_BITS'd1981790147, `RNS_PRIME_BITS'd1869463650, `RNS_PRIME_BITS'd1134712329, `RNS_PRIME_BITS'd617071312, `RNS_PRIME_BITS'd1082506074, `RNS_PRIME_BITS'd868206324, `RNS_PRIME_BITS'd741081945, `RNS_PRIME_BITS'd584967224},
			'{`RNS_PRIME_BITS'd77, `RNS_PRIME_BITS'd764311327, `RNS_PRIME_BITS'd1879454363, `RNS_PRIME_BITS'd451097162, `RNS_PRIME_BITS'd963259320, `RNS_PRIME_BITS'd883302316, `RNS_PRIME_BITS'd1915298618, `RNS_PRIME_BITS'd1072701021, `RNS_PRIME_BITS'd338373351, `RNS_PRIME_BITS'd1136416059, `RNS_PRIME_BITS'd1690878566},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd1759625170, `RNS_PRIME_BITS'd1907931650, `RNS_PRIME_BITS'd477155584, `RNS_PRIME_BITS'd1074539447, `RNS_PRIME_BITS'd1806492734, `RNS_PRIME_BITS'd1298771737, `RNS_PRIME_BITS'd742830755, `RNS_PRIME_BITS'd233432035, `RNS_PRIME_BITS'd1488325428, `RNS_PRIME_BITS'd1797028726},
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd110176105, `RNS_PRIME_BITS'd474987895, `RNS_PRIME_BITS'd1741901560, `RNS_PRIME_BITS'd1192334265, `RNS_PRIME_BITS'd255604877, `RNS_PRIME_BITS'd1963120340, `RNS_PRIME_BITS'd116073025, `RNS_PRIME_BITS'd354982278, `RNS_PRIME_BITS'd1687350507, `RNS_PRIME_BITS'd1615971935},
			'{`RNS_PRIME_BITS'd102, `RNS_PRIME_BITS'd547524178, `RNS_PRIME_BITS'd1230455148, `RNS_PRIME_BITS'd324594532, `RNS_PRIME_BITS'd956658810, `RNS_PRIME_BITS'd1997861131, `RNS_PRIME_BITS'd322249427, `RNS_PRIME_BITS'd1424582828, `RNS_PRIME_BITS'd576947822, `RNS_PRIME_BITS'd2041780307, `RNS_PRIME_BITS'd531051162},
			'{`RNS_PRIME_BITS'd19, `RNS_PRIME_BITS'd1755326225, `RNS_PRIME_BITS'd2059248419, `RNS_PRIME_BITS'd599236922, `RNS_PRIME_BITS'd305270234, `RNS_PRIME_BITS'd801251863, `RNS_PRIME_BITS'd525642616, `RNS_PRIME_BITS'd1014348323, `RNS_PRIME_BITS'd1560772533, `RNS_PRIME_BITS'd2042093837, `RNS_PRIME_BITS'd1679968384},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd1117054723, `RNS_PRIME_BITS'd392965232, `RNS_PRIME_BITS'd1661708401, `RNS_PRIME_BITS'd733484050, `RNS_PRIME_BITS'd873389187, `RNS_PRIME_BITS'd1822674099, `RNS_PRIME_BITS'd595934223, `RNS_PRIME_BITS'd1100991334, `RNS_PRIME_BITS'd2000006977, `RNS_PRIME_BITS'd164282191},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd873415029, `RNS_PRIME_BITS'd1416757354, `RNS_PRIME_BITS'd2119451090, `RNS_PRIME_BITS'd1530627789, `RNS_PRIME_BITS'd1234759544, `RNS_PRIME_BITS'd970702151, `RNS_PRIME_BITS'd1383551822, `RNS_PRIME_BITS'd608699265, `RNS_PRIME_BITS'd2025803221, `RNS_PRIME_BITS'd1030775517},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd355109779, `RNS_PRIME_BITS'd1944773438, `RNS_PRIME_BITS'd1641807579, `RNS_PRIME_BITS'd40722566, `RNS_PRIME_BITS'd1790487069, `RNS_PRIME_BITS'd1265712404, `RNS_PRIME_BITS'd695811555, `RNS_PRIME_BITS'd364584294, `RNS_PRIME_BITS'd1338027655, `RNS_PRIME_BITS'd1503978156},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd1330285964, `RNS_PRIME_BITS'd245082899, `RNS_PRIME_BITS'd333460392, `RNS_PRIME_BITS'd551160321, `RNS_PRIME_BITS'd136615721, `RNS_PRIME_BITS'd1407638400, `RNS_PRIME_BITS'd1545525455, `RNS_PRIME_BITS'd2062451649, `RNS_PRIME_BITS'd1934837338, `RNS_PRIME_BITS'd116329066},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd901459116, `RNS_PRIME_BITS'd1147981710, `RNS_PRIME_BITS'd1776034545, `RNS_PRIME_BITS'd1565239439, `RNS_PRIME_BITS'd1945133948, `RNS_PRIME_BITS'd762952382, `RNS_PRIME_BITS'd34623499, `RNS_PRIME_BITS'd2117469183, `RNS_PRIME_BITS'd590977683, `RNS_PRIME_BITS'd149686646},
			'{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd42624479, `RNS_PRIME_BITS'd967227428, `RNS_PRIME_BITS'd1425081841, `RNS_PRIME_BITS'd514154763, `RNS_PRIME_BITS'd554991597, `RNS_PRIME_BITS'd2128623742, `RNS_PRIME_BITS'd2106811745, `RNS_PRIME_BITS'd924078218, `RNS_PRIME_BITS'd1077757630, `RNS_PRIME_BITS'd1538491376},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd961583221, `RNS_PRIME_BITS'd1485558273, `RNS_PRIME_BITS'd249086558, `RNS_PRIME_BITS'd918072858, `RNS_PRIME_BITS'd1295268023, `RNS_PRIME_BITS'd1582475445, `RNS_PRIME_BITS'd767877127, `RNS_PRIME_BITS'd1850075585, `RNS_PRIME_BITS'd2074078634, `RNS_PRIME_BITS'd1115595790},
			'{`RNS_PRIME_BITS'd28, `RNS_PRIME_BITS'd2032672218, `RNS_PRIME_BITS'd115955423, `RNS_PRIME_BITS'd1763196099, `RNS_PRIME_BITS'd807542637, `RNS_PRIME_BITS'd1207250116, `RNS_PRIME_BITS'd2016593392, `RNS_PRIME_BITS'd659126444, `RNS_PRIME_BITS'd2057148765, `RNS_PRIME_BITS'd1901774972, `RNS_PRIME_BITS'd1353141292},
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd1660953538, `RNS_PRIME_BITS'd585552958, `RNS_PRIME_BITS'd242272109, `RNS_PRIME_BITS'd1992321453, `RNS_PRIME_BITS'd2053877646, `RNS_PRIME_BITS'd1589753902, `RNS_PRIME_BITS'd2045206131, `RNS_PRIME_BITS'd980478047, `RNS_PRIME_BITS'd1220771174, `RNS_PRIME_BITS'd357242888},
			'{`RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd1264194384, `RNS_PRIME_BITS'd1080633195, `RNS_PRIME_BITS'd206011688, `RNS_PRIME_BITS'd2029509785, `RNS_PRIME_BITS'd83910918, `RNS_PRIME_BITS'd418285876, `RNS_PRIME_BITS'd1233675354, `RNS_PRIME_BITS'd507058184, `RNS_PRIME_BITS'd1943734012, `RNS_PRIME_BITS'd1895479845},
			'{`RNS_PRIME_BITS'd219, `RNS_PRIME_BITS'd1960653297, `RNS_PRIME_BITS'd1443782123, `RNS_PRIME_BITS'd1904197865, `RNS_PRIME_BITS'd1829024041, `RNS_PRIME_BITS'd489780005, `RNS_PRIME_BITS'd1440461339, `RNS_PRIME_BITS'd1395544982, `RNS_PRIME_BITS'd182931571, `RNS_PRIME_BITS'd886670302, `RNS_PRIME_BITS'd1657905200},
			'{`RNS_PRIME_BITS'd27, `RNS_PRIME_BITS'd615456589, `RNS_PRIME_BITS'd400978795, `RNS_PRIME_BITS'd1672506762, `RNS_PRIME_BITS'd1707738, `RNS_PRIME_BITS'd1624010767, `RNS_PRIME_BITS'd1608587393, `RNS_PRIME_BITS'd1813940954, `RNS_PRIME_BITS'd1327923721, `RNS_PRIME_BITS'd310644219, `RNS_PRIME_BITS'd163236766},
			'{`RNS_PRIME_BITS'd213, `RNS_PRIME_BITS'd44420466, `RNS_PRIME_BITS'd1585811054, `RNS_PRIME_BITS'd1390728917, `RNS_PRIME_BITS'd1345185166, `RNS_PRIME_BITS'd275417299, `RNS_PRIME_BITS'd632397777, `RNS_PRIME_BITS'd1222865969, `RNS_PRIME_BITS'd1689931663, `RNS_PRIME_BITS'd1016353521, `RNS_PRIME_BITS'd743618593},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd1611326066, `RNS_PRIME_BITS'd354506087, `RNS_PRIME_BITS'd2004096401, `RNS_PRIME_BITS'd1162217418, `RNS_PRIME_BITS'd1722057271, `RNS_PRIME_BITS'd798189785, `RNS_PRIME_BITS'd1106392084, `RNS_PRIME_BITS'd539777139, `RNS_PRIME_BITS'd1930188078, `RNS_PRIME_BITS'd171939123},
			'{`RNS_PRIME_BITS'd54, `RNS_PRIME_BITS'd656575985, `RNS_PRIME_BITS'd1025116930, `RNS_PRIME_BITS'd845173269, `RNS_PRIME_BITS'd2137754810, `RNS_PRIME_BITS'd953052890, `RNS_PRIME_BITS'd1265755320, `RNS_PRIME_BITS'd175856921, `RNS_PRIME_BITS'd1285635300, `RNS_PRIME_BITS'd370744456, `RNS_PRIME_BITS'd155225031},
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd1499545593, `RNS_PRIME_BITS'd1698398402, `RNS_PRIME_BITS'd1968289269, `RNS_PRIME_BITS'd394990771, `RNS_PRIME_BITS'd634543754, `RNS_PRIME_BITS'd1788527753, `RNS_PRIME_BITS'd77650491, `RNS_PRIME_BITS'd669713681, `RNS_PRIME_BITS'd482748218, `RNS_PRIME_BITS'd927892699},
			'{`RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd1116676029, `RNS_PRIME_BITS'd1504639209, `RNS_PRIME_BITS'd1161739390, `RNS_PRIME_BITS'd229159739, `RNS_PRIME_BITS'd1081953270, `RNS_PRIME_BITS'd462419066, `RNS_PRIME_BITS'd1858799108, `RNS_PRIME_BITS'd17356827, `RNS_PRIME_BITS'd658169400, `RNS_PRIME_BITS'd1996101824},
			'{`RNS_PRIME_BITS'd177, `RNS_PRIME_BITS'd1813744972, `RNS_PRIME_BITS'd1972979682, `RNS_PRIME_BITS'd206865569, `RNS_PRIME_BITS'd451041711, `RNS_PRIME_BITS'd393958967, `RNS_PRIME_BITS'd1093636343, `RNS_PRIME_BITS'd913354707, `RNS_PRIME_BITS'd1027265014, `RNS_PRIME_BITS'd175440921, `RNS_PRIME_BITS'd829915829},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd396645382, `RNS_PRIME_BITS'd1791657634, `RNS_PRIME_BITS'd1413541989, `RNS_PRIME_BITS'd2081875639, `RNS_PRIME_BITS'd794161257, `RNS_PRIME_BITS'd1270258990, `RNS_PRIME_BITS'd516680554, `RNS_PRIME_BITS'd669076203, `RNS_PRIME_BITS'd421308264, `RNS_PRIME_BITS'd1086822439},
			'{`RNS_PRIME_BITS'd83, `RNS_PRIME_BITS'd69134841, `RNS_PRIME_BITS'd1821416425, `RNS_PRIME_BITS'd50752640, `RNS_PRIME_BITS'd1655191859, `RNS_PRIME_BITS'd1921993674, `RNS_PRIME_BITS'd451196014, `RNS_PRIME_BITS'd1000662686, `RNS_PRIME_BITS'd647048807, `RNS_PRIME_BITS'd932182495, `RNS_PRIME_BITS'd391797855},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd877304277, `RNS_PRIME_BITS'd159977213, `RNS_PRIME_BITS'd290077813, `RNS_PRIME_BITS'd1810063376, `RNS_PRIME_BITS'd566748967, `RNS_PRIME_BITS'd639538435, `RNS_PRIME_BITS'd1484063037, `RNS_PRIME_BITS'd55792857, `RNS_PRIME_BITS'd1714473259, `RNS_PRIME_BITS'd2144012390},
			'{`RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd50571811, `RNS_PRIME_BITS'd2115181952, `RNS_PRIME_BITS'd562019831, `RNS_PRIME_BITS'd1154612085, `RNS_PRIME_BITS'd1786639521, `RNS_PRIME_BITS'd1925769136, `RNS_PRIME_BITS'd1728369768, `RNS_PRIME_BITS'd2085135257, `RNS_PRIME_BITS'd295310129, `RNS_PRIME_BITS'd1336425779},
			'{`RNS_PRIME_BITS'd115, `RNS_PRIME_BITS'd4002933, `RNS_PRIME_BITS'd2075292787, `RNS_PRIME_BITS'd1983768083, `RNS_PRIME_BITS'd1023350667, `RNS_PRIME_BITS'd176309237, `RNS_PRIME_BITS'd1593277516, `RNS_PRIME_BITS'd1382104874, `RNS_PRIME_BITS'd1523915141, `RNS_PRIME_BITS'd848075412, `RNS_PRIME_BITS'd765646662},
			'{`RNS_PRIME_BITS'd94, `RNS_PRIME_BITS'd573597879, `RNS_PRIME_BITS'd1344174270, `RNS_PRIME_BITS'd2100132974, `RNS_PRIME_BITS'd777005688, `RNS_PRIME_BITS'd574185762, `RNS_PRIME_BITS'd131328332, `RNS_PRIME_BITS'd1169773623, `RNS_PRIME_BITS'd887851340, `RNS_PRIME_BITS'd1125787949, `RNS_PRIME_BITS'd353599546},
			'{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd59147011, `RNS_PRIME_BITS'd2123418675, `RNS_PRIME_BITS'd435046516, `RNS_PRIME_BITS'd88645780, `RNS_PRIME_BITS'd260032417, `RNS_PRIME_BITS'd2104091640, `RNS_PRIME_BITS'd1823306947, `RNS_PRIME_BITS'd2109457066, `RNS_PRIME_BITS'd1163737865, `RNS_PRIME_BITS'd1767353290},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd1394136953, `RNS_PRIME_BITS'd1173090837, `RNS_PRIME_BITS'd995824257, `RNS_PRIME_BITS'd437515366, `RNS_PRIME_BITS'd1208997909, `RNS_PRIME_BITS'd822456584, `RNS_PRIME_BITS'd1874625716, `RNS_PRIME_BITS'd1431298095, `RNS_PRIME_BITS'd1665451287, `RNS_PRIME_BITS'd1553222695},
			'{`RNS_PRIME_BITS'd149, `RNS_PRIME_BITS'd941632951, `RNS_PRIME_BITS'd1694944408, `RNS_PRIME_BITS'd1546038111, `RNS_PRIME_BITS'd524895673, `RNS_PRIME_BITS'd1239252466, `RNS_PRIME_BITS'd90055778, `RNS_PRIME_BITS'd731280767, `RNS_PRIME_BITS'd600741851, `RNS_PRIME_BITS'd1738927365, `RNS_PRIME_BITS'd1588148031},
			'{`RNS_PRIME_BITS'd140, `RNS_PRIME_BITS'd2140093298, `RNS_PRIME_BITS'd759046863, `RNS_PRIME_BITS'd264915896, `RNS_PRIME_BITS'd1772042254, `RNS_PRIME_BITS'd1259854095, `RNS_PRIME_BITS'd1802742692, `RNS_PRIME_BITS'd61004180, `RNS_PRIME_BITS'd242090628, `RNS_PRIME_BITS'd1451307179, `RNS_PRIME_BITS'd943837035},
			'{`RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd1542577651, `RNS_PRIME_BITS'd1685711514, `RNS_PRIME_BITS'd2039463678, `RNS_PRIME_BITS'd1047434922, `RNS_PRIME_BITS'd978140117, `RNS_PRIME_BITS'd1472757042, `RNS_PRIME_BITS'd399486371, `RNS_PRIME_BITS'd736407238, `RNS_PRIME_BITS'd364857629, `RNS_PRIME_BITS'd1254229217},
			'{`RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd1137828556, `RNS_PRIME_BITS'd113535793, `RNS_PRIME_BITS'd1693338984, `RNS_PRIME_BITS'd1238765823, `RNS_PRIME_BITS'd842844032, `RNS_PRIME_BITS'd515131391, `RNS_PRIME_BITS'd484363258, `RNS_PRIME_BITS'd1716973785, `RNS_PRIME_BITS'd1293120823, `RNS_PRIME_BITS'd841842457},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd1942253647, `RNS_PRIME_BITS'd1409329318, `RNS_PRIME_BITS'd46804831, `RNS_PRIME_BITS'd42942124, `RNS_PRIME_BITS'd1636484991, `RNS_PRIME_BITS'd2018352455, `RNS_PRIME_BITS'd1294487706, `RNS_PRIME_BITS'd998147012, `RNS_PRIME_BITS'd1586352206, `RNS_PRIME_BITS'd993498128},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1594438390, `RNS_PRIME_BITS'd1080892916, `RNS_PRIME_BITS'd557127875, `RNS_PRIME_BITS'd242313701, `RNS_PRIME_BITS'd1211072570, `RNS_PRIME_BITS'd486053531, `RNS_PRIME_BITS'd1201661802, `RNS_PRIME_BITS'd594106034, `RNS_PRIME_BITS'd1655116100, `RNS_PRIME_BITS'd1950842557},
			'{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd2147313512, `RNS_PRIME_BITS'd1755989622, `RNS_PRIME_BITS'd1345883903, `RNS_PRIME_BITS'd1367395951, `RNS_PRIME_BITS'd1649356752, `RNS_PRIME_BITS'd704887596, `RNS_PRIME_BITS'd1802515947, `RNS_PRIME_BITS'd1069986885, `RNS_PRIME_BITS'd1221222533, `RNS_PRIME_BITS'd600509576},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd1817052548, `RNS_PRIME_BITS'd2094546834, `RNS_PRIME_BITS'd669268230, `RNS_PRIME_BITS'd1903185293, `RNS_PRIME_BITS'd2109203059, `RNS_PRIME_BITS'd1709674595, `RNS_PRIME_BITS'd915795313, `RNS_PRIME_BITS'd806329581, `RNS_PRIME_BITS'd40649261, `RNS_PRIME_BITS'd606640892},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd1991277784, `RNS_PRIME_BITS'd1310508345, `RNS_PRIME_BITS'd194811738, `RNS_PRIME_BITS'd1427910660, `RNS_PRIME_BITS'd35507526, `RNS_PRIME_BITS'd640823705, `RNS_PRIME_BITS'd1190738917, `RNS_PRIME_BITS'd367925886, `RNS_PRIME_BITS'd1474154399, `RNS_PRIME_BITS'd1976764288},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd782812247, `RNS_PRIME_BITS'd2005003043, `RNS_PRIME_BITS'd1309802650, `RNS_PRIME_BITS'd996789255, `RNS_PRIME_BITS'd1034092333, `RNS_PRIME_BITS'd1772860827, `RNS_PRIME_BITS'd1000786930, `RNS_PRIME_BITS'd123268731, `RNS_PRIME_BITS'd1192478917, `RNS_PRIME_BITS'd560204155},
			'{`RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd135906172, `RNS_PRIME_BITS'd1412319986, `RNS_PRIME_BITS'd1948097938, `RNS_PRIME_BITS'd1710814283, `RNS_PRIME_BITS'd928823477, `RNS_PRIME_BITS'd389121690, `RNS_PRIME_BITS'd1779430027, `RNS_PRIME_BITS'd1901937128, `RNS_PRIME_BITS'd370311231, `RNS_PRIME_BITS'd1214189046},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd841038518, `RNS_PRIME_BITS'd289672111, `RNS_PRIME_BITS'd375180356, `RNS_PRIME_BITS'd1567343535, `RNS_PRIME_BITS'd23853187, `RNS_PRIME_BITS'd915960474, `RNS_PRIME_BITS'd240489248, `RNS_PRIME_BITS'd1539865624, `RNS_PRIME_BITS'd1618503395, `RNS_PRIME_BITS'd1659823052}
		},
		'{
			'{`RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd2110550228, `RNS_PRIME_BITS'd1722149111, `RNS_PRIME_BITS'd999667849, `RNS_PRIME_BITS'd532899428, `RNS_PRIME_BITS'd1553179927, `RNS_PRIME_BITS'd2040290224, `RNS_PRIME_BITS'd975561682, `RNS_PRIME_BITS'd1830870858, `RNS_PRIME_BITS'd1873700450, `RNS_PRIME_BITS'd1910852744},
			'{`RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd2129301944, `RNS_PRIME_BITS'd1638985049, `RNS_PRIME_BITS'd1615408981, `RNS_PRIME_BITS'd753080299, `RNS_PRIME_BITS'd701719901, `RNS_PRIME_BITS'd1502899173, `RNS_PRIME_BITS'd898913524, `RNS_PRIME_BITS'd274828075, `RNS_PRIME_BITS'd210409048, `RNS_PRIME_BITS'd1032426123},
			'{`RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd1143708976, `RNS_PRIME_BITS'd978579843, `RNS_PRIME_BITS'd839923132, `RNS_PRIME_BITS'd845293986, `RNS_PRIME_BITS'd26339099, `RNS_PRIME_BITS'd1832545566, `RNS_PRIME_BITS'd1972569442, `RNS_PRIME_BITS'd564907987, `RNS_PRIME_BITS'd974858260, `RNS_PRIME_BITS'd507515759},
			'{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd1838882159, `RNS_PRIME_BITS'd76011792, `RNS_PRIME_BITS'd1569607090, `RNS_PRIME_BITS'd742879251, `RNS_PRIME_BITS'd1750380170, `RNS_PRIME_BITS'd2010053405, `RNS_PRIME_BITS'd265545663, `RNS_PRIME_BITS'd1017354991, `RNS_PRIME_BITS'd1524533295, `RNS_PRIME_BITS'd716204455},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd2105298764, `RNS_PRIME_BITS'd1471580670, `RNS_PRIME_BITS'd2003231283, `RNS_PRIME_BITS'd1044022036, `RNS_PRIME_BITS'd348752518, `RNS_PRIME_BITS'd698417353, `RNS_PRIME_BITS'd1500535600, `RNS_PRIME_BITS'd965423605, `RNS_PRIME_BITS'd1915012469, `RNS_PRIME_BITS'd1996709144},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd619801035, `RNS_PRIME_BITS'd782007668, `RNS_PRIME_BITS'd816887802, `RNS_PRIME_BITS'd849822566, `RNS_PRIME_BITS'd739448663, `RNS_PRIME_BITS'd1443722027, `RNS_PRIME_BITS'd389041925, `RNS_PRIME_BITS'd651329317, `RNS_PRIME_BITS'd1328400050, `RNS_PRIME_BITS'd309827063},
			'{`RNS_PRIME_BITS'd206, `RNS_PRIME_BITS'd794681083, `RNS_PRIME_BITS'd1758671978, `RNS_PRIME_BITS'd388829693, `RNS_PRIME_BITS'd987961512, `RNS_PRIME_BITS'd888591969, `RNS_PRIME_BITS'd610031167, `RNS_PRIME_BITS'd1365164089, `RNS_PRIME_BITS'd978360583, `RNS_PRIME_BITS'd2129970825, `RNS_PRIME_BITS'd765190713},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1328671547, `RNS_PRIME_BITS'd246824953, `RNS_PRIME_BITS'd431275491, `RNS_PRIME_BITS'd605765246, `RNS_PRIME_BITS'd693368348, `RNS_PRIME_BITS'd1477659904, `RNS_PRIME_BITS'd2146336963, `RNS_PRIME_BITS'd1359400799, `RNS_PRIME_BITS'd1937009915, `RNS_PRIME_BITS'd927522827},
			'{`RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd57406560, `RNS_PRIME_BITS'd582533808, `RNS_PRIME_BITS'd130814149, `RNS_PRIME_BITS'd567980090, `RNS_PRIME_BITS'd1569800392, `RNS_PRIME_BITS'd679132985, `RNS_PRIME_BITS'd303044825, `RNS_PRIME_BITS'd1509142993, `RNS_PRIME_BITS'd159647058, `RNS_PRIME_BITS'd1958980030},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd438618986, `RNS_PRIME_BITS'd2124186313, `RNS_PRIME_BITS'd254016143, `RNS_PRIME_BITS'd524235090, `RNS_PRIME_BITS'd1112755321, `RNS_PRIME_BITS'd774025118, `RNS_PRIME_BITS'd2071933749, `RNS_PRIME_BITS'd244853563, `RNS_PRIME_BITS'd102873346, `RNS_PRIME_BITS'd914169442},
			'{`RNS_PRIME_BITS'd152, `RNS_PRIME_BITS'd1172837580, `RNS_PRIME_BITS'd1017828612, `RNS_PRIME_BITS'd660584570, `RNS_PRIME_BITS'd467401747, `RNS_PRIME_BITS'd1219012245, `RNS_PRIME_BITS'd675137241, `RNS_PRIME_BITS'd142410138, `RNS_PRIME_BITS'd2122234197, `RNS_PRIME_BITS'd601489443, `RNS_PRIME_BITS'd988969898},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd695648387, `RNS_PRIME_BITS'd1274590505, `RNS_PRIME_BITS'd600982728, `RNS_PRIME_BITS'd433103425, `RNS_PRIME_BITS'd2016123870, `RNS_PRIME_BITS'd692035776, `RNS_PRIME_BITS'd2082713122, `RNS_PRIME_BITS'd177892363, `RNS_PRIME_BITS'd671824567, `RNS_PRIME_BITS'd236309105},
			'{`RNS_PRIME_BITS'd174, `RNS_PRIME_BITS'd604330433, `RNS_PRIME_BITS'd2035929063, `RNS_PRIME_BITS'd1506445507, `RNS_PRIME_BITS'd528747556, `RNS_PRIME_BITS'd475091879, `RNS_PRIME_BITS'd2029890290, `RNS_PRIME_BITS'd788239302, `RNS_PRIME_BITS'd1831066174, `RNS_PRIME_BITS'd1249974132, `RNS_PRIME_BITS'd1714038324},
			'{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd2019189855, `RNS_PRIME_BITS'd1714454654, `RNS_PRIME_BITS'd579355062, `RNS_PRIME_BITS'd1587946537, `RNS_PRIME_BITS'd1066762236, `RNS_PRIME_BITS'd325808629, `RNS_PRIME_BITS'd575109967, `RNS_PRIME_BITS'd926022203, `RNS_PRIME_BITS'd1030352876, `RNS_PRIME_BITS'd1759968861},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd1738680099, `RNS_PRIME_BITS'd649757504, `RNS_PRIME_BITS'd2087811899, `RNS_PRIME_BITS'd1247466235, `RNS_PRIME_BITS'd1555607486, `RNS_PRIME_BITS'd1548661104, `RNS_PRIME_BITS'd1818734790, `RNS_PRIME_BITS'd191730041, `RNS_PRIME_BITS'd17892876, `RNS_PRIME_BITS'd606316738},
			'{`RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd870023649, `RNS_PRIME_BITS'd1119466787, `RNS_PRIME_BITS'd1196822847, `RNS_PRIME_BITS'd1307591471, `RNS_PRIME_BITS'd702006335, `RNS_PRIME_BITS'd1980439017, `RNS_PRIME_BITS'd824700098, `RNS_PRIME_BITS'd1091404214, `RNS_PRIME_BITS'd1794617198, `RNS_PRIME_BITS'd1201435568},
			'{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd481387912, `RNS_PRIME_BITS'd1006538441, `RNS_PRIME_BITS'd1837970192, `RNS_PRIME_BITS'd12108181, `RNS_PRIME_BITS'd1083969199, `RNS_PRIME_BITS'd985153668, `RNS_PRIME_BITS'd257107127, `RNS_PRIME_BITS'd1816446847, `RNS_PRIME_BITS'd162743922, `RNS_PRIME_BITS'd1939746247},
			'{`RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd757528441, `RNS_PRIME_BITS'd803544833, `RNS_PRIME_BITS'd123300694, `RNS_PRIME_BITS'd643469593, `RNS_PRIME_BITS'd670756904, `RNS_PRIME_BITS'd381908047, `RNS_PRIME_BITS'd42133797, `RNS_PRIME_BITS'd1533690942, `RNS_PRIME_BITS'd646057027, `RNS_PRIME_BITS'd1084451174},
			'{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd1665060078, `RNS_PRIME_BITS'd15051646, `RNS_PRIME_BITS'd1793722621, `RNS_PRIME_BITS'd1546974591, `RNS_PRIME_BITS'd617071047, `RNS_PRIME_BITS'd556067091, `RNS_PRIME_BITS'd1011444201, `RNS_PRIME_BITS'd1612142892, `RNS_PRIME_BITS'd1369615129, `RNS_PRIME_BITS'd1371056440},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd564071341, `RNS_PRIME_BITS'd1750744336, `RNS_PRIME_BITS'd487883017, `RNS_PRIME_BITS'd986036689, `RNS_PRIME_BITS'd1230493654, `RNS_PRIME_BITS'd443095192, `RNS_PRIME_BITS'd595179459, `RNS_PRIME_BITS'd1913402093, `RNS_PRIME_BITS'd1079425714, `RNS_PRIME_BITS'd62539456},
			'{`RNS_PRIME_BITS'd161, `RNS_PRIME_BITS'd797650456, `RNS_PRIME_BITS'd819800400, `RNS_PRIME_BITS'd149563950, `RNS_PRIME_BITS'd1017311971, `RNS_PRIME_BITS'd828195520, `RNS_PRIME_BITS'd243231637, `RNS_PRIME_BITS'd1594182033, `RNS_PRIME_BITS'd1325352760, `RNS_PRIME_BITS'd2108643044, `RNS_PRIME_BITS'd188218960},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd566665698, `RNS_PRIME_BITS'd995999548, `RNS_PRIME_BITS'd1436223500, `RNS_PRIME_BITS'd1071821487, `RNS_PRIME_BITS'd1626062709, `RNS_PRIME_BITS'd1190171477, `RNS_PRIME_BITS'd1192192635, `RNS_PRIME_BITS'd1041633442, `RNS_PRIME_BITS'd1356208944, `RNS_PRIME_BITS'd1595292078},
			'{`RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd1069538846, `RNS_PRIME_BITS'd1440479555, `RNS_PRIME_BITS'd964094715, `RNS_PRIME_BITS'd2015419361, `RNS_PRIME_BITS'd926676223, `RNS_PRIME_BITS'd837491928, `RNS_PRIME_BITS'd1538656458, `RNS_PRIME_BITS'd2007342038, `RNS_PRIME_BITS'd2014624705, `RNS_PRIME_BITS'd863620233},
			'{`RNS_PRIME_BITS'd32, `RNS_PRIME_BITS'd1872969846, `RNS_PRIME_BITS'd1405607800, `RNS_PRIME_BITS'd357424905, `RNS_PRIME_BITS'd559851995, `RNS_PRIME_BITS'd1766244905, `RNS_PRIME_BITS'd606445012, `RNS_PRIME_BITS'd705023616, `RNS_PRIME_BITS'd698481148, `RNS_PRIME_BITS'd2120132974, `RNS_PRIME_BITS'd1879753738},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd990994856, `RNS_PRIME_BITS'd1350825992, `RNS_PRIME_BITS'd660408957, `RNS_PRIME_BITS'd1524214037, `RNS_PRIME_BITS'd1045734136, `RNS_PRIME_BITS'd1802988279, `RNS_PRIME_BITS'd726129993, `RNS_PRIME_BITS'd93963335, `RNS_PRIME_BITS'd188563254, `RNS_PRIME_BITS'd543878303},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd1966812310, `RNS_PRIME_BITS'd2056360637, `RNS_PRIME_BITS'd897057228, `RNS_PRIME_BITS'd487668072, `RNS_PRIME_BITS'd1849571421, `RNS_PRIME_BITS'd838761593, `RNS_PRIME_BITS'd1908809754, `RNS_PRIME_BITS'd426238081, `RNS_PRIME_BITS'd1705600854, `RNS_PRIME_BITS'd1929780323},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd249827822, `RNS_PRIME_BITS'd2063055506, `RNS_PRIME_BITS'd903330376, `RNS_PRIME_BITS'd1985575130, `RNS_PRIME_BITS'd622435062, `RNS_PRIME_BITS'd550662787, `RNS_PRIME_BITS'd1256385395, `RNS_PRIME_BITS'd2119957118, `RNS_PRIME_BITS'd1178256475, `RNS_PRIME_BITS'd52020526},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd726515733, `RNS_PRIME_BITS'd604779166, `RNS_PRIME_BITS'd1480718190, `RNS_PRIME_BITS'd1833355609, `RNS_PRIME_BITS'd2053843334, `RNS_PRIME_BITS'd382827394, `RNS_PRIME_BITS'd1888093051, `RNS_PRIME_BITS'd282767684, `RNS_PRIME_BITS'd1417586066, `RNS_PRIME_BITS'd908868540},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd1190074285, `RNS_PRIME_BITS'd329912932, `RNS_PRIME_BITS'd1495580858, `RNS_PRIME_BITS'd2127810203, `RNS_PRIME_BITS'd563072674, `RNS_PRIME_BITS'd1579414323, `RNS_PRIME_BITS'd733765447, `RNS_PRIME_BITS'd247891300, `RNS_PRIME_BITS'd918434589, `RNS_PRIME_BITS'd1631077461},
			'{`RNS_PRIME_BITS'd250, `RNS_PRIME_BITS'd657737713, `RNS_PRIME_BITS'd418756999, `RNS_PRIME_BITS'd669241465, `RNS_PRIME_BITS'd1342048858, `RNS_PRIME_BITS'd103369633, `RNS_PRIME_BITS'd1363556183, `RNS_PRIME_BITS'd768679511, `RNS_PRIME_BITS'd283180663, `RNS_PRIME_BITS'd1081354292, `RNS_PRIME_BITS'd1414651605},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd368330405, `RNS_PRIME_BITS'd1022220406, `RNS_PRIME_BITS'd954509746, `RNS_PRIME_BITS'd973726281, `RNS_PRIME_BITS'd1203697433, `RNS_PRIME_BITS'd2049241416, `RNS_PRIME_BITS'd440447715, `RNS_PRIME_BITS'd400712242, `RNS_PRIME_BITS'd1898274856, `RNS_PRIME_BITS'd1392674349},
			'{`RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd1419673164, `RNS_PRIME_BITS'd1480022475, `RNS_PRIME_BITS'd1703685595, `RNS_PRIME_BITS'd184244689, `RNS_PRIME_BITS'd2102134578, `RNS_PRIME_BITS'd2109641780, `RNS_PRIME_BITS'd824531322, `RNS_PRIME_BITS'd1440640937, `RNS_PRIME_BITS'd92209613, `RNS_PRIME_BITS'd162313921},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd604245432, `RNS_PRIME_BITS'd491162767, `RNS_PRIME_BITS'd235268169, `RNS_PRIME_BITS'd1244217216, `RNS_PRIME_BITS'd900342339, `RNS_PRIME_BITS'd429128151, `RNS_PRIME_BITS'd982261016, `RNS_PRIME_BITS'd1635454096, `RNS_PRIME_BITS'd577369776, `RNS_PRIME_BITS'd447700181},
			'{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd419073016, `RNS_PRIME_BITS'd1813862106, `RNS_PRIME_BITS'd1257894537, `RNS_PRIME_BITS'd397211051, `RNS_PRIME_BITS'd1428040779, `RNS_PRIME_BITS'd2095377683, `RNS_PRIME_BITS'd864629636, `RNS_PRIME_BITS'd1208147894, `RNS_PRIME_BITS'd1232823458, `RNS_PRIME_BITS'd1562312453},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd1428971954, `RNS_PRIME_BITS'd1867767814, `RNS_PRIME_BITS'd530385897, `RNS_PRIME_BITS'd894398625, `RNS_PRIME_BITS'd1809846362, `RNS_PRIME_BITS'd137438335, `RNS_PRIME_BITS'd99895886, `RNS_PRIME_BITS'd423019830, `RNS_PRIME_BITS'd303127306, `RNS_PRIME_BITS'd1470692548},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd1687614984, `RNS_PRIME_BITS'd709280857, `RNS_PRIME_BITS'd1342532931, `RNS_PRIME_BITS'd1760527589, `RNS_PRIME_BITS'd1148164666, `RNS_PRIME_BITS'd769204672, `RNS_PRIME_BITS'd220924129, `RNS_PRIME_BITS'd601999986, `RNS_PRIME_BITS'd1897487815, `RNS_PRIME_BITS'd2068509710},
			'{`RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd954409419, `RNS_PRIME_BITS'd1757057320, `RNS_PRIME_BITS'd1144645785, `RNS_PRIME_BITS'd548145161, `RNS_PRIME_BITS'd1646514035, `RNS_PRIME_BITS'd412508002, `RNS_PRIME_BITS'd1966156222, `RNS_PRIME_BITS'd422465534, `RNS_PRIME_BITS'd78725657, `RNS_PRIME_BITS'd1222910613},
			'{`RNS_PRIME_BITS'd74, `RNS_PRIME_BITS'd1399847152, `RNS_PRIME_BITS'd1833287656, `RNS_PRIME_BITS'd1327366429, `RNS_PRIME_BITS'd645878241, `RNS_PRIME_BITS'd1695769720, `RNS_PRIME_BITS'd783334765, `RNS_PRIME_BITS'd2093798455, `RNS_PRIME_BITS'd1798031938, `RNS_PRIME_BITS'd359261796, `RNS_PRIME_BITS'd580828799},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd1212695587, `RNS_PRIME_BITS'd1484801920, `RNS_PRIME_BITS'd1498757522, `RNS_PRIME_BITS'd840450833, `RNS_PRIME_BITS'd737118709, `RNS_PRIME_BITS'd1656945872, `RNS_PRIME_BITS'd1748329974, `RNS_PRIME_BITS'd1744500512, `RNS_PRIME_BITS'd2119548962, `RNS_PRIME_BITS'd1636409584},
			'{`RNS_PRIME_BITS'd202, `RNS_PRIME_BITS'd1290309463, `RNS_PRIME_BITS'd1972942824, `RNS_PRIME_BITS'd2010044655, `RNS_PRIME_BITS'd682674352, `RNS_PRIME_BITS'd53708544, `RNS_PRIME_BITS'd1688718488, `RNS_PRIME_BITS'd2099854708, `RNS_PRIME_BITS'd591650138, `RNS_PRIME_BITS'd1821345941, `RNS_PRIME_BITS'd1248012241},
			'{`RNS_PRIME_BITS'd233, `RNS_PRIME_BITS'd131710303, `RNS_PRIME_BITS'd1993987715, `RNS_PRIME_BITS'd2051282882, `RNS_PRIME_BITS'd45333268, `RNS_PRIME_BITS'd302970267, `RNS_PRIME_BITS'd1058537647, `RNS_PRIME_BITS'd1070212953, `RNS_PRIME_BITS'd1086596263, `RNS_PRIME_BITS'd1185669667, `RNS_PRIME_BITS'd554513430},
			'{`RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd1501786709, `RNS_PRIME_BITS'd1869109985, `RNS_PRIME_BITS'd202914531, `RNS_PRIME_BITS'd1895453977, `RNS_PRIME_BITS'd742527237, `RNS_PRIME_BITS'd1635039913, `RNS_PRIME_BITS'd1576296687, `RNS_PRIME_BITS'd1638648932, `RNS_PRIME_BITS'd1600889350, `RNS_PRIME_BITS'd1759384411},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd999273190, `RNS_PRIME_BITS'd2070844445, `RNS_PRIME_BITS'd861050475, `RNS_PRIME_BITS'd1491712965, `RNS_PRIME_BITS'd813221858, `RNS_PRIME_BITS'd984867860, `RNS_PRIME_BITS'd1653260604, `RNS_PRIME_BITS'd878801800, `RNS_PRIME_BITS'd879540287, `RNS_PRIME_BITS'd191450223},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd532550233, `RNS_PRIME_BITS'd1327897855, `RNS_PRIME_BITS'd1279008922, `RNS_PRIME_BITS'd2048128415, `RNS_PRIME_BITS'd1888260297, `RNS_PRIME_BITS'd989651243, `RNS_PRIME_BITS'd1870423980, `RNS_PRIME_BITS'd1448459171, `RNS_PRIME_BITS'd1209167554, `RNS_PRIME_BITS'd1352078228},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1237750355, `RNS_PRIME_BITS'd191612023, `RNS_PRIME_BITS'd65447791, `RNS_PRIME_BITS'd318336440, `RNS_PRIME_BITS'd797044206, `RNS_PRIME_BITS'd1834998783, `RNS_PRIME_BITS'd1079056222, `RNS_PRIME_BITS'd1305317978, `RNS_PRIME_BITS'd758318031, `RNS_PRIME_BITS'd344740188},
			'{`RNS_PRIME_BITS'd192, `RNS_PRIME_BITS'd170463767, `RNS_PRIME_BITS'd1724044163, `RNS_PRIME_BITS'd1501965744, `RNS_PRIME_BITS'd820165498, `RNS_PRIME_BITS'd1011304463, `RNS_PRIME_BITS'd2119886881, `RNS_PRIME_BITS'd325527626, `RNS_PRIME_BITS'd752574849, `RNS_PRIME_BITS'd1465412733, `RNS_PRIME_BITS'd1283396089},
			'{`RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd793607665, `RNS_PRIME_BITS'd1988776824, `RNS_PRIME_BITS'd1242107079, `RNS_PRIME_BITS'd527540060, `RNS_PRIME_BITS'd72035215, `RNS_PRIME_BITS'd1695453503, `RNS_PRIME_BITS'd1842827729, `RNS_PRIME_BITS'd468629171, `RNS_PRIME_BITS'd728734694, `RNS_PRIME_BITS'd1276129449},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd1798961482, `RNS_PRIME_BITS'd1739969704, `RNS_PRIME_BITS'd1501560594, `RNS_PRIME_BITS'd1287542248, `RNS_PRIME_BITS'd684419942, `RNS_PRIME_BITS'd1018855866, `RNS_PRIME_BITS'd1615131826, `RNS_PRIME_BITS'd66308458, `RNS_PRIME_BITS'd260569056, `RNS_PRIME_BITS'd290522827},
			'{`RNS_PRIME_BITS'd130, `RNS_PRIME_BITS'd927449603, `RNS_PRIME_BITS'd1875728858, `RNS_PRIME_BITS'd1177411113, `RNS_PRIME_BITS'd1003048664, `RNS_PRIME_BITS'd1578315522, `RNS_PRIME_BITS'd1696532957, `RNS_PRIME_BITS'd1905910587, `RNS_PRIME_BITS'd74099818, `RNS_PRIME_BITS'd1572443018, `RNS_PRIME_BITS'd1220132623},
			'{`RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd1293203516, `RNS_PRIME_BITS'd172846845, `RNS_PRIME_BITS'd1207637146, `RNS_PRIME_BITS'd186595044, `RNS_PRIME_BITS'd239335674, `RNS_PRIME_BITS'd1066718425, `RNS_PRIME_BITS'd410038680, `RNS_PRIME_BITS'd1739338584, `RNS_PRIME_BITS'd985552131, `RNS_PRIME_BITS'd39270801},
			'{`RNS_PRIME_BITS'd155, `RNS_PRIME_BITS'd1376067929, `RNS_PRIME_BITS'd1537808658, `RNS_PRIME_BITS'd1597482381, `RNS_PRIME_BITS'd1252224832, `RNS_PRIME_BITS'd1815597825, `RNS_PRIME_BITS'd1359306658, `RNS_PRIME_BITS'd1691889137, `RNS_PRIME_BITS'd1606150984, `RNS_PRIME_BITS'd546458997, `RNS_PRIME_BITS'd1230626089},
			'{`RNS_PRIME_BITS'd75, `RNS_PRIME_BITS'd294592480, `RNS_PRIME_BITS'd68254058, `RNS_PRIME_BITS'd2045572413, `RNS_PRIME_BITS'd1582726490, `RNS_PRIME_BITS'd806139582, `RNS_PRIME_BITS'd1790592449, `RNS_PRIME_BITS'd760220325, `RNS_PRIME_BITS'd200986787, `RNS_PRIME_BITS'd1014529300, `RNS_PRIME_BITS'd1944773851},
			'{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd156088985, `RNS_PRIME_BITS'd95500170, `RNS_PRIME_BITS'd1908908193, `RNS_PRIME_BITS'd1229775075, `RNS_PRIME_BITS'd573774165, `RNS_PRIME_BITS'd635759498, `RNS_PRIME_BITS'd395900530, `RNS_PRIME_BITS'd1306598371, `RNS_PRIME_BITS'd194780596, `RNS_PRIME_BITS'd1320225974},
			'{`RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd1497148278, `RNS_PRIME_BITS'd186556355, `RNS_PRIME_BITS'd955712373, `RNS_PRIME_BITS'd1996296427, `RNS_PRIME_BITS'd1025720640, `RNS_PRIME_BITS'd1444815208, `RNS_PRIME_BITS'd270420625, `RNS_PRIME_BITS'd899456512, `RNS_PRIME_BITS'd349886599, `RNS_PRIME_BITS'd676720427},
			'{`RNS_PRIME_BITS'd97, `RNS_PRIME_BITS'd1306471650, `RNS_PRIME_BITS'd2022829342, `RNS_PRIME_BITS'd1456015930, `RNS_PRIME_BITS'd1865431418, `RNS_PRIME_BITS'd1481574512, `RNS_PRIME_BITS'd109864796, `RNS_PRIME_BITS'd1342375658, `RNS_PRIME_BITS'd1589255329, `RNS_PRIME_BITS'd1255472078, `RNS_PRIME_BITS'd1362139157},
			'{`RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd505970387, `RNS_PRIME_BITS'd1356884376, `RNS_PRIME_BITS'd1545487606, `RNS_PRIME_BITS'd293127918, `RNS_PRIME_BITS'd669906709, `RNS_PRIME_BITS'd293293168, `RNS_PRIME_BITS'd795985671, `RNS_PRIME_BITS'd15527131, `RNS_PRIME_BITS'd113694653, `RNS_PRIME_BITS'd451445947},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd949150133, `RNS_PRIME_BITS'd120972581, `RNS_PRIME_BITS'd1791213139, `RNS_PRIME_BITS'd1801245249, `RNS_PRIME_BITS'd1701022176, `RNS_PRIME_BITS'd737608443, `RNS_PRIME_BITS'd1466471468, `RNS_PRIME_BITS'd929238933, `RNS_PRIME_BITS'd1308679709, `RNS_PRIME_BITS'd1843083092},
			'{`RNS_PRIME_BITS'd216, `RNS_PRIME_BITS'd1065038128, `RNS_PRIME_BITS'd97158433, `RNS_PRIME_BITS'd1114028516, `RNS_PRIME_BITS'd699701463, `RNS_PRIME_BITS'd2050390163, `RNS_PRIME_BITS'd1962005329, `RNS_PRIME_BITS'd1187652640, `RNS_PRIME_BITS'd1904240392, `RNS_PRIME_BITS'd1663468063, `RNS_PRIME_BITS'd1801841561},
			'{`RNS_PRIME_BITS'd232, `RNS_PRIME_BITS'd2037385759, `RNS_PRIME_BITS'd1765111518, `RNS_PRIME_BITS'd54005447, `RNS_PRIME_BITS'd766495802, `RNS_PRIME_BITS'd715250119, `RNS_PRIME_BITS'd1653804360, `RNS_PRIME_BITS'd1474602261, `RNS_PRIME_BITS'd74240402, `RNS_PRIME_BITS'd447783940, `RNS_PRIME_BITS'd1211073467},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd547690395, `RNS_PRIME_BITS'd1045363286, `RNS_PRIME_BITS'd1032220652, `RNS_PRIME_BITS'd920248116, `RNS_PRIME_BITS'd1828804801, `RNS_PRIME_BITS'd1038813682, `RNS_PRIME_BITS'd762294407, `RNS_PRIME_BITS'd452132682, `RNS_PRIME_BITS'd1731110774, `RNS_PRIME_BITS'd720752137},
			'{`RNS_PRIME_BITS'd20, `RNS_PRIME_BITS'd1515018158, `RNS_PRIME_BITS'd1253039887, `RNS_PRIME_BITS'd18958806, `RNS_PRIME_BITS'd1709378496, `RNS_PRIME_BITS'd93787655, `RNS_PRIME_BITS'd978495501, `RNS_PRIME_BITS'd905468019, `RNS_PRIME_BITS'd9988371, `RNS_PRIME_BITS'd96294344, `RNS_PRIME_BITS'd1233998733},
			'{`RNS_PRIME_BITS'd247, `RNS_PRIME_BITS'd1254420141, `RNS_PRIME_BITS'd378301072, `RNS_PRIME_BITS'd71925555, `RNS_PRIME_BITS'd884367919, `RNS_PRIME_BITS'd213832555, `RNS_PRIME_BITS'd326805075, `RNS_PRIME_BITS'd785328188, `RNS_PRIME_BITS'd1430454074, `RNS_PRIME_BITS'd1088223894, `RNS_PRIME_BITS'd1206129988},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd603187420, `RNS_PRIME_BITS'd940312975, `RNS_PRIME_BITS'd632137340, `RNS_PRIME_BITS'd1396065490, `RNS_PRIME_BITS'd1300358994, `RNS_PRIME_BITS'd973137737, `RNS_PRIME_BITS'd1843866585, `RNS_PRIME_BITS'd1310423022, `RNS_PRIME_BITS'd1119212180, `RNS_PRIME_BITS'd68292664},
			'{`RNS_PRIME_BITS'd238, `RNS_PRIME_BITS'd1530324037, `RNS_PRIME_BITS'd100112297, `RNS_PRIME_BITS'd787258385, `RNS_PRIME_BITS'd1168747153, `RNS_PRIME_BITS'd1696397126, `RNS_PRIME_BITS'd1037497317, `RNS_PRIME_BITS'd1208919114, `RNS_PRIME_BITS'd1295060874, `RNS_PRIME_BITS'd1836223655, `RNS_PRIME_BITS'd47663904}
		}
	},
	'{
		'{
			'{`RNS_PRIME_BITS'd31, `RNS_PRIME_BITS'd194696075, `RNS_PRIME_BITS'd2060302498, `RNS_PRIME_BITS'd82728389, `RNS_PRIME_BITS'd439200745, `RNS_PRIME_BITS'd199167574, `RNS_PRIME_BITS'd1018979385, `RNS_PRIME_BITS'd444259819, `RNS_PRIME_BITS'd816792377, `RNS_PRIME_BITS'd35859490, `RNS_PRIME_BITS'd737695627},
			'{`RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd374351703, `RNS_PRIME_BITS'd1696495122, `RNS_PRIME_BITS'd1700399344, `RNS_PRIME_BITS'd970227529, `RNS_PRIME_BITS'd1468121814, `RNS_PRIME_BITS'd1322752092, `RNS_PRIME_BITS'd649280504, `RNS_PRIME_BITS'd1240606164, `RNS_PRIME_BITS'd1404704941, `RNS_PRIME_BITS'd242632142},
			'{`RNS_PRIME_BITS'd229, `RNS_PRIME_BITS'd1989607565, `RNS_PRIME_BITS'd1719251453, `RNS_PRIME_BITS'd90539947, `RNS_PRIME_BITS'd1441524485, `RNS_PRIME_BITS'd1695395048, `RNS_PRIME_BITS'd1942129095, `RNS_PRIME_BITS'd822970348, `RNS_PRIME_BITS'd1481551325, `RNS_PRIME_BITS'd823884731, `RNS_PRIME_BITS'd1659015304},
			'{`RNS_PRIME_BITS'd145, `RNS_PRIME_BITS'd1213485156, `RNS_PRIME_BITS'd724534082, `RNS_PRIME_BITS'd612290505, `RNS_PRIME_BITS'd483430963, `RNS_PRIME_BITS'd1514986211, `RNS_PRIME_BITS'd989890522, `RNS_PRIME_BITS'd1596450073, `RNS_PRIME_BITS'd912103023, `RNS_PRIME_BITS'd42584731, `RNS_PRIME_BITS'd565249089},
			'{`RNS_PRIME_BITS'd47, `RNS_PRIME_BITS'd1174086677, `RNS_PRIME_BITS'd1755044050, `RNS_PRIME_BITS'd1294260305, `RNS_PRIME_BITS'd497364496, `RNS_PRIME_BITS'd866272432, `RNS_PRIME_BITS'd2037553853, `RNS_PRIME_BITS'd782477094, `RNS_PRIME_BITS'd424803860, `RNS_PRIME_BITS'd1422242550, `RNS_PRIME_BITS'd1025817260},
			'{`RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd1735917560, `RNS_PRIME_BITS'd712008187, `RNS_PRIME_BITS'd237483994, `RNS_PRIME_BITS'd1448655249, `RNS_PRIME_BITS'd1050035780, `RNS_PRIME_BITS'd332802255, `RNS_PRIME_BITS'd1060344472, `RNS_PRIME_BITS'd1618657303, `RNS_PRIME_BITS'd1801709110, `RNS_PRIME_BITS'd360727220},
			'{`RNS_PRIME_BITS'd219, `RNS_PRIME_BITS'd801237025, `RNS_PRIME_BITS'd2050167408, `RNS_PRIME_BITS'd308909792, `RNS_PRIME_BITS'd1395232827, `RNS_PRIME_BITS'd543207486, `RNS_PRIME_BITS'd1853730580, `RNS_PRIME_BITS'd1991829268, `RNS_PRIME_BITS'd688173292, `RNS_PRIME_BITS'd2034707373, `RNS_PRIME_BITS'd1681213823},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd470305790, `RNS_PRIME_BITS'd1782975752, `RNS_PRIME_BITS'd729460484, `RNS_PRIME_BITS'd1068726870, `RNS_PRIME_BITS'd1349396655, `RNS_PRIME_BITS'd1508428172, `RNS_PRIME_BITS'd1200206602, `RNS_PRIME_BITS'd821039318, `RNS_PRIME_BITS'd45681605, `RNS_PRIME_BITS'd953333869},
			'{`RNS_PRIME_BITS'd201, `RNS_PRIME_BITS'd1689558788, `RNS_PRIME_BITS'd1519594416, `RNS_PRIME_BITS'd47347478, `RNS_PRIME_BITS'd1997332060, `RNS_PRIME_BITS'd35835091, `RNS_PRIME_BITS'd741568614, `RNS_PRIME_BITS'd140709962, `RNS_PRIME_BITS'd779046918, `RNS_PRIME_BITS'd826137934, `RNS_PRIME_BITS'd1428573171},
			'{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1238876179, `RNS_PRIME_BITS'd861747159, `RNS_PRIME_BITS'd1882256500, `RNS_PRIME_BITS'd1854447557, `RNS_PRIME_BITS'd33067001, `RNS_PRIME_BITS'd2045767491, `RNS_PRIME_BITS'd2023095682, `RNS_PRIME_BITS'd669812059, `RNS_PRIME_BITS'd1032129870, `RNS_PRIME_BITS'd2703558},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd1445056051, `RNS_PRIME_BITS'd871429424, `RNS_PRIME_BITS'd1103190308, `RNS_PRIME_BITS'd1823746342, `RNS_PRIME_BITS'd882751157, `RNS_PRIME_BITS'd1012202940, `RNS_PRIME_BITS'd341027723, `RNS_PRIME_BITS'd1644004709, `RNS_PRIME_BITS'd2024023420, `RNS_PRIME_BITS'd1568722053},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd6384100, `RNS_PRIME_BITS'd941190001, `RNS_PRIME_BITS'd1940466509, `RNS_PRIME_BITS'd100497516, `RNS_PRIME_BITS'd1104355284, `RNS_PRIME_BITS'd1790033930, `RNS_PRIME_BITS'd686119614, `RNS_PRIME_BITS'd1940635540, `RNS_PRIME_BITS'd1203262265, `RNS_PRIME_BITS'd35892535},
			'{`RNS_PRIME_BITS'd220, `RNS_PRIME_BITS'd1168350968, `RNS_PRIME_BITS'd507243856, `RNS_PRIME_BITS'd2021993277, `RNS_PRIME_BITS'd1886991642, `RNS_PRIME_BITS'd1279894373, `RNS_PRIME_BITS'd135403194, `RNS_PRIME_BITS'd195815254, `RNS_PRIME_BITS'd1383318536, `RNS_PRIME_BITS'd1702381996, `RNS_PRIME_BITS'd1618534321},
			'{`RNS_PRIME_BITS'd86, `RNS_PRIME_BITS'd612116218, `RNS_PRIME_BITS'd447499598, `RNS_PRIME_BITS'd309566020, `RNS_PRIME_BITS'd1568904359, `RNS_PRIME_BITS'd221724701, `RNS_PRIME_BITS'd90871238, `RNS_PRIME_BITS'd1316400403, `RNS_PRIME_BITS'd673801197, `RNS_PRIME_BITS'd134353639, `RNS_PRIME_BITS'd821400007},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd122083856, `RNS_PRIME_BITS'd951061445, `RNS_PRIME_BITS'd1908640337, `RNS_PRIME_BITS'd1029126052, `RNS_PRIME_BITS'd222300657, `RNS_PRIME_BITS'd1456499969, `RNS_PRIME_BITS'd1427415160, `RNS_PRIME_BITS'd474281196, `RNS_PRIME_BITS'd875473710, `RNS_PRIME_BITS'd535360449},
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd366060953, `RNS_PRIME_BITS'd203523950, `RNS_PRIME_BITS'd1317674688, `RNS_PRIME_BITS'd1487412974, `RNS_PRIME_BITS'd780568852, `RNS_PRIME_BITS'd12189015, `RNS_PRIME_BITS'd120525056, `RNS_PRIME_BITS'd448825163, `RNS_PRIME_BITS'd1243803783, `RNS_PRIME_BITS'd171410388},
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd831438452, `RNS_PRIME_BITS'd246732979, `RNS_PRIME_BITS'd699219664, `RNS_PRIME_BITS'd1773281056, `RNS_PRIME_BITS'd638427284, `RNS_PRIME_BITS'd41054675, `RNS_PRIME_BITS'd185757691, `RNS_PRIME_BITS'd1979332317, `RNS_PRIME_BITS'd86672268, `RNS_PRIME_BITS'd1457305023},
			'{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd1561641664, `RNS_PRIME_BITS'd1378076090, `RNS_PRIME_BITS'd546654075, `RNS_PRIME_BITS'd1399958391, `RNS_PRIME_BITS'd893979190, `RNS_PRIME_BITS'd883764098, `RNS_PRIME_BITS'd939546168, `RNS_PRIME_BITS'd331359640, `RNS_PRIME_BITS'd2109759261, `RNS_PRIME_BITS'd808305431},
			'{`RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd759618172, `RNS_PRIME_BITS'd1323692621, `RNS_PRIME_BITS'd641500902, `RNS_PRIME_BITS'd1349043972, `RNS_PRIME_BITS'd2087107446, `RNS_PRIME_BITS'd1583567685, `RNS_PRIME_BITS'd81417488, `RNS_PRIME_BITS'd1273566470, `RNS_PRIME_BITS'd2036560478, `RNS_PRIME_BITS'd1015891554},
			'{`RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd720073991, `RNS_PRIME_BITS'd2033751660, `RNS_PRIME_BITS'd419483890, `RNS_PRIME_BITS'd828778002, `RNS_PRIME_BITS'd1177680023, `RNS_PRIME_BITS'd1061660784, `RNS_PRIME_BITS'd1190788793, `RNS_PRIME_BITS'd1251325708, `RNS_PRIME_BITS'd1998013280, `RNS_PRIME_BITS'd1116897775},
			'{`RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd1356916561, `RNS_PRIME_BITS'd873438397, `RNS_PRIME_BITS'd722043381, `RNS_PRIME_BITS'd960812949, `RNS_PRIME_BITS'd587907123, `RNS_PRIME_BITS'd1845173464, `RNS_PRIME_BITS'd178844159, `RNS_PRIME_BITS'd556005356, `RNS_PRIME_BITS'd730577106, `RNS_PRIME_BITS'd602881725},
			'{`RNS_PRIME_BITS'd90, `RNS_PRIME_BITS'd908656677, `RNS_PRIME_BITS'd150043102, `RNS_PRIME_BITS'd1365393962, `RNS_PRIME_BITS'd2054985161, `RNS_PRIME_BITS'd1279062800, `RNS_PRIME_BITS'd1929027214, `RNS_PRIME_BITS'd1635240377, `RNS_PRIME_BITS'd825677997, `RNS_PRIME_BITS'd1266062834, `RNS_PRIME_BITS'd1974290835},
			'{`RNS_PRIME_BITS'd126, `RNS_PRIME_BITS'd1712662486, `RNS_PRIME_BITS'd1292575444, `RNS_PRIME_BITS'd1118508252, `RNS_PRIME_BITS'd1990860009, `RNS_PRIME_BITS'd914661085, `RNS_PRIME_BITS'd1548824054, `RNS_PRIME_BITS'd43384459, `RNS_PRIME_BITS'd158324149, `RNS_PRIME_BITS'd1618209596, `RNS_PRIME_BITS'd1694142340},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd1117284082, `RNS_PRIME_BITS'd2053272228, `RNS_PRIME_BITS'd1644010299, `RNS_PRIME_BITS'd662777964, `RNS_PRIME_BITS'd2054118730, `RNS_PRIME_BITS'd1752314571, `RNS_PRIME_BITS'd989955561, `RNS_PRIME_BITS'd1387821852, `RNS_PRIME_BITS'd1366490698, `RNS_PRIME_BITS'd1076385929},
			'{`RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd1863191856, `RNS_PRIME_BITS'd103003952, `RNS_PRIME_BITS'd1775533903, `RNS_PRIME_BITS'd2038757092, `RNS_PRIME_BITS'd1904182858, `RNS_PRIME_BITS'd1515559419, `RNS_PRIME_BITS'd992898587, `RNS_PRIME_BITS'd1201662396, `RNS_PRIME_BITS'd1229549280, `RNS_PRIME_BITS'd1162705990},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd1533981961, `RNS_PRIME_BITS'd2025706356, `RNS_PRIME_BITS'd1715379271, `RNS_PRIME_BITS'd769786813, `RNS_PRIME_BITS'd500561489, `RNS_PRIME_BITS'd1842904497, `RNS_PRIME_BITS'd1845987112, `RNS_PRIME_BITS'd2144467332, `RNS_PRIME_BITS'd1554294293, `RNS_PRIME_BITS'd2098442982},
			'{`RNS_PRIME_BITS'd56, `RNS_PRIME_BITS'd1533174716, `RNS_PRIME_BITS'd1317351157, `RNS_PRIME_BITS'd2055365765, `RNS_PRIME_BITS'd1494002858, `RNS_PRIME_BITS'd1815205203, `RNS_PRIME_BITS'd1174159037, `RNS_PRIME_BITS'd1595079530, `RNS_PRIME_BITS'd121893430, `RNS_PRIME_BITS'd82865862, `RNS_PRIME_BITS'd70495657},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1177975178, `RNS_PRIME_BITS'd1783454984, `RNS_PRIME_BITS'd2147020409, `RNS_PRIME_BITS'd344232922, `RNS_PRIME_BITS'd1471651844, `RNS_PRIME_BITS'd1018907210, `RNS_PRIME_BITS'd1320243887, `RNS_PRIME_BITS'd810430885, `RNS_PRIME_BITS'd1539177095, `RNS_PRIME_BITS'd1531727760},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd1179715763, `RNS_PRIME_BITS'd1659069973, `RNS_PRIME_BITS'd229998048, `RNS_PRIME_BITS'd79500857, `RNS_PRIME_BITS'd1033265161, `RNS_PRIME_BITS'd2128544231, `RNS_PRIME_BITS'd1924445104, `RNS_PRIME_BITS'd1286502494, `RNS_PRIME_BITS'd103248575, `RNS_PRIME_BITS'd969861422},
			'{`RNS_PRIME_BITS'd3, `RNS_PRIME_BITS'd1529199458, `RNS_PRIME_BITS'd1134865089, `RNS_PRIME_BITS'd1138755299, `RNS_PRIME_BITS'd1749738016, `RNS_PRIME_BITS'd1347111703, `RNS_PRIME_BITS'd856731473, `RNS_PRIME_BITS'd1366434580, `RNS_PRIME_BITS'd555068228, `RNS_PRIME_BITS'd1273645171, `RNS_PRIME_BITS'd451643648},
			'{`RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd2027264733, `RNS_PRIME_BITS'd2017570980, `RNS_PRIME_BITS'd401575901, `RNS_PRIME_BITS'd530148286, `RNS_PRIME_BITS'd186617009, `RNS_PRIME_BITS'd2024954824, `RNS_PRIME_BITS'd213349046, `RNS_PRIME_BITS'd1648926136, `RNS_PRIME_BITS'd1022384850, `RNS_PRIME_BITS'd198834507},
			'{`RNS_PRIME_BITS'd69, `RNS_PRIME_BITS'd997453221, `RNS_PRIME_BITS'd1284561451, `RNS_PRIME_BITS'd616152262, `RNS_PRIME_BITS'd1149278255, `RNS_PRIME_BITS'd676575321, `RNS_PRIME_BITS'd1329872757, `RNS_PRIME_BITS'd1261303829, `RNS_PRIME_BITS'd716041462, `RNS_PRIME_BITS'd1531466762, `RNS_PRIME_BITS'd916968946},
			'{`RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd1456154083, `RNS_PRIME_BITS'd1345121295, `RNS_PRIME_BITS'd1009073918, `RNS_PRIME_BITS'd886896888, `RNS_PRIME_BITS'd1636768070, `RNS_PRIME_BITS'd2014615209, `RNS_PRIME_BITS'd968402202, `RNS_PRIME_BITS'd2089023679, `RNS_PRIME_BITS'd87676709, `RNS_PRIME_BITS'd1305602516},
			'{`RNS_PRIME_BITS'd164, `RNS_PRIME_BITS'd1408161112, `RNS_PRIME_BITS'd1674502898, `RNS_PRIME_BITS'd365146251, `RNS_PRIME_BITS'd20115630, `RNS_PRIME_BITS'd406288528, `RNS_PRIME_BITS'd1912823087, `RNS_PRIME_BITS'd108939319, `RNS_PRIME_BITS'd425059557, `RNS_PRIME_BITS'd2025694180, `RNS_PRIME_BITS'd1164995614},
			'{`RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd1813126663, `RNS_PRIME_BITS'd1237681120, `RNS_PRIME_BITS'd1750139962, `RNS_PRIME_BITS'd802189914, `RNS_PRIME_BITS'd760938321, `RNS_PRIME_BITS'd1129864153, `RNS_PRIME_BITS'd666023594, `RNS_PRIME_BITS'd1231732887, `RNS_PRIME_BITS'd907691071, `RNS_PRIME_BITS'd1216922722},
			'{`RNS_PRIME_BITS'd224, `RNS_PRIME_BITS'd1132073771, `RNS_PRIME_BITS'd620146647, `RNS_PRIME_BITS'd1782999443, `RNS_PRIME_BITS'd1803748509, `RNS_PRIME_BITS'd568728513, `RNS_PRIME_BITS'd2039322147, `RNS_PRIME_BITS'd2012683352, `RNS_PRIME_BITS'd1551049847, `RNS_PRIME_BITS'd1272775921, `RNS_PRIME_BITS'd791327078},
			'{`RNS_PRIME_BITS'd212, `RNS_PRIME_BITS'd1620225369, `RNS_PRIME_BITS'd856725124, `RNS_PRIME_BITS'd849267490, `RNS_PRIME_BITS'd1863139568, `RNS_PRIME_BITS'd1394147207, `RNS_PRIME_BITS'd1784577441, `RNS_PRIME_BITS'd2037024441, `RNS_PRIME_BITS'd1362800672, `RNS_PRIME_BITS'd1177047477, `RNS_PRIME_BITS'd1846577282},
			'{`RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd793579694, `RNS_PRIME_BITS'd1527001438, `RNS_PRIME_BITS'd2011963482, `RNS_PRIME_BITS'd1946075888, `RNS_PRIME_BITS'd1425374308, `RNS_PRIME_BITS'd1579522935, `RNS_PRIME_BITS'd204798715, `RNS_PRIME_BITS'd233328130, `RNS_PRIME_BITS'd1897063024, `RNS_PRIME_BITS'd1532253084},
			'{`RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd639728460, `RNS_PRIME_BITS'd1868470216, `RNS_PRIME_BITS'd527671976, `RNS_PRIME_BITS'd2002444714, `RNS_PRIME_BITS'd1175263851, `RNS_PRIME_BITS'd1928363754, `RNS_PRIME_BITS'd1222403150, `RNS_PRIME_BITS'd578904461, `RNS_PRIME_BITS'd1211311735, `RNS_PRIME_BITS'd504488370},
			'{`RNS_PRIME_BITS'd237, `RNS_PRIME_BITS'd1396198292, `RNS_PRIME_BITS'd1920590771, `RNS_PRIME_BITS'd387776744, `RNS_PRIME_BITS'd963163635, `RNS_PRIME_BITS'd1203233787, `RNS_PRIME_BITS'd1484894886, `RNS_PRIME_BITS'd1502544141, `RNS_PRIME_BITS'd104204490, `RNS_PRIME_BITS'd1362839063, `RNS_PRIME_BITS'd1844052458},
			'{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd485420777, `RNS_PRIME_BITS'd807501472, `RNS_PRIME_BITS'd1757068898, `RNS_PRIME_BITS'd1358003415, `RNS_PRIME_BITS'd1675687172, `RNS_PRIME_BITS'd662827380, `RNS_PRIME_BITS'd1915528076, `RNS_PRIME_BITS'd1757954929, `RNS_PRIME_BITS'd1405633615, `RNS_PRIME_BITS'd1116677626},
			'{`RNS_PRIME_BITS'd19, `RNS_PRIME_BITS'd1015946329, `RNS_PRIME_BITS'd1019987263, `RNS_PRIME_BITS'd1174476985, `RNS_PRIME_BITS'd1885452558, `RNS_PRIME_BITS'd1725297415, `RNS_PRIME_BITS'd1229007112, `RNS_PRIME_BITS'd111014336, `RNS_PRIME_BITS'd1373728089, `RNS_PRIME_BITS'd998561906, `RNS_PRIME_BITS'd1841410565},
			'{`RNS_PRIME_BITS'd243, `RNS_PRIME_BITS'd659763983, `RNS_PRIME_BITS'd5902460, `RNS_PRIME_BITS'd359945354, `RNS_PRIME_BITS'd999155403, `RNS_PRIME_BITS'd1823605536, `RNS_PRIME_BITS'd301313136, `RNS_PRIME_BITS'd1537588749, `RNS_PRIME_BITS'd2130633339, `RNS_PRIME_BITS'd451643617, `RNS_PRIME_BITS'd1842199681},
			'{`RNS_PRIME_BITS'd245, `RNS_PRIME_BITS'd577637347, `RNS_PRIME_BITS'd1359947184, `RNS_PRIME_BITS'd1328518975, `RNS_PRIME_BITS'd1455650682, `RNS_PRIME_BITS'd1992552230, `RNS_PRIME_BITS'd1748513462, `RNS_PRIME_BITS'd91281715, `RNS_PRIME_BITS'd634139283, `RNS_PRIME_BITS'd1087718144, `RNS_PRIME_BITS'd1401902809},
			'{`RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd1661032155, `RNS_PRIME_BITS'd500810373, `RNS_PRIME_BITS'd1636512422, `RNS_PRIME_BITS'd175021434, `RNS_PRIME_BITS'd1802461381, `RNS_PRIME_BITS'd1579381933, `RNS_PRIME_BITS'd132456626, `RNS_PRIME_BITS'd337340874, `RNS_PRIME_BITS'd103598397, `RNS_PRIME_BITS'd140787404},
			'{`RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd1630985590, `RNS_PRIME_BITS'd672875555, `RNS_PRIME_BITS'd1783753433, `RNS_PRIME_BITS'd1014947771, `RNS_PRIME_BITS'd526414536, `RNS_PRIME_BITS'd1850696922, `RNS_PRIME_BITS'd824229110, `RNS_PRIME_BITS'd1360378682, `RNS_PRIME_BITS'd618593197, `RNS_PRIME_BITS'd364243142},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd1723690242, `RNS_PRIME_BITS'd469996204, `RNS_PRIME_BITS'd2057066390, `RNS_PRIME_BITS'd826778132, `RNS_PRIME_BITS'd1806048511, `RNS_PRIME_BITS'd500184242, `RNS_PRIME_BITS'd965058738, `RNS_PRIME_BITS'd1511343746, `RNS_PRIME_BITS'd1616960181, `RNS_PRIME_BITS'd427464610},
			'{`RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd2090431652, `RNS_PRIME_BITS'd949564075, `RNS_PRIME_BITS'd96121591, `RNS_PRIME_BITS'd919343373, `RNS_PRIME_BITS'd1907509843, `RNS_PRIME_BITS'd1953384801, `RNS_PRIME_BITS'd1457490910, `RNS_PRIME_BITS'd478934848, `RNS_PRIME_BITS'd2116550331, `RNS_PRIME_BITS'd879990775},
			'{`RNS_PRIME_BITS'd45, `RNS_PRIME_BITS'd68594092, `RNS_PRIME_BITS'd1950774255, `RNS_PRIME_BITS'd698674139, `RNS_PRIME_BITS'd822634792, `RNS_PRIME_BITS'd1758999004, `RNS_PRIME_BITS'd1264923480, `RNS_PRIME_BITS'd1356561501, `RNS_PRIME_BITS'd1516568707, `RNS_PRIME_BITS'd1242380800, `RNS_PRIME_BITS'd1051566862},
			'{`RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd276244453, `RNS_PRIME_BITS'd1223269848, `RNS_PRIME_BITS'd222604456, `RNS_PRIME_BITS'd1210366788, `RNS_PRIME_BITS'd899044363, `RNS_PRIME_BITS'd1018288932, `RNS_PRIME_BITS'd78485193, `RNS_PRIME_BITS'd1389010213, `RNS_PRIME_BITS'd848347554, `RNS_PRIME_BITS'd1414453716},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd254312299, `RNS_PRIME_BITS'd1535482010, `RNS_PRIME_BITS'd527451978, `RNS_PRIME_BITS'd95004208, `RNS_PRIME_BITS'd1585445351, `RNS_PRIME_BITS'd1272346785, `RNS_PRIME_BITS'd483004783, `RNS_PRIME_BITS'd321164175, `RNS_PRIME_BITS'd97063170, `RNS_PRIME_BITS'd1219460139},
			'{`RNS_PRIME_BITS'd80, `RNS_PRIME_BITS'd1905216912, `RNS_PRIME_BITS'd159693917, `RNS_PRIME_BITS'd76681201, `RNS_PRIME_BITS'd245429092, `RNS_PRIME_BITS'd1174836922, `RNS_PRIME_BITS'd1252805571, `RNS_PRIME_BITS'd276449714, `RNS_PRIME_BITS'd888504768, `RNS_PRIME_BITS'd1489064321, `RNS_PRIME_BITS'd380049315},
			'{`RNS_PRIME_BITS'd32, `RNS_PRIME_BITS'd2142312425, `RNS_PRIME_BITS'd1569865949, `RNS_PRIME_BITS'd974250149, `RNS_PRIME_BITS'd1754951921, `RNS_PRIME_BITS'd1116129849, `RNS_PRIME_BITS'd1477098398, `RNS_PRIME_BITS'd626451913, `RNS_PRIME_BITS'd1736848206, `RNS_PRIME_BITS'd549050356, `RNS_PRIME_BITS'd341514572},
			'{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1307339339, `RNS_PRIME_BITS'd1200318051, `RNS_PRIME_BITS'd1135547408, `RNS_PRIME_BITS'd324721317, `RNS_PRIME_BITS'd695034078, `RNS_PRIME_BITS'd1149126389, `RNS_PRIME_BITS'd1685944029, `RNS_PRIME_BITS'd419228638, `RNS_PRIME_BITS'd1805059831, `RNS_PRIME_BITS'd294425532},
			'{`RNS_PRIME_BITS'd175, `RNS_PRIME_BITS'd1301817278, `RNS_PRIME_BITS'd1107521354, `RNS_PRIME_BITS'd1376702860, `RNS_PRIME_BITS'd1792726430, `RNS_PRIME_BITS'd204189914, `RNS_PRIME_BITS'd149799757, `RNS_PRIME_BITS'd588941338, `RNS_PRIME_BITS'd114641712, `RNS_PRIME_BITS'd1363985959, `RNS_PRIME_BITS'd155727161},
			'{`RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd1453088379, `RNS_PRIME_BITS'd254768500, `RNS_PRIME_BITS'd925610389, `RNS_PRIME_BITS'd1719573924, `RNS_PRIME_BITS'd967382750, `RNS_PRIME_BITS'd1122238909, `RNS_PRIME_BITS'd989059247, `RNS_PRIME_BITS'd2000687997, `RNS_PRIME_BITS'd1417628163, `RNS_PRIME_BITS'd1816330104},
			'{`RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd1038095229, `RNS_PRIME_BITS'd1818413900, `RNS_PRIME_BITS'd1814275570, `RNS_PRIME_BITS'd1743932620, `RNS_PRIME_BITS'd1647149675, `RNS_PRIME_BITS'd951137760, `RNS_PRIME_BITS'd903984566, `RNS_PRIME_BITS'd1950044445, `RNS_PRIME_BITS'd1214769201, `RNS_PRIME_BITS'd1163177753},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd551165231, `RNS_PRIME_BITS'd424409902, `RNS_PRIME_BITS'd1989305716, `RNS_PRIME_BITS'd1122450322, `RNS_PRIME_BITS'd95144970, `RNS_PRIME_BITS'd2090439576, `RNS_PRIME_BITS'd1314627921, `RNS_PRIME_BITS'd31945130, `RNS_PRIME_BITS'd1185254040, `RNS_PRIME_BITS'd2077622591},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd632554148, `RNS_PRIME_BITS'd1580330817, `RNS_PRIME_BITS'd1937666267, `RNS_PRIME_BITS'd1878109348, `RNS_PRIME_BITS'd1700580858, `RNS_PRIME_BITS'd2132459452, `RNS_PRIME_BITS'd423792449, `RNS_PRIME_BITS'd1246328674, `RNS_PRIME_BITS'd544758867, `RNS_PRIME_BITS'd1045449225},
			'{`RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd1555160323, `RNS_PRIME_BITS'd473196449, `RNS_PRIME_BITS'd257488132, `RNS_PRIME_BITS'd1413736043, `RNS_PRIME_BITS'd604628799, `RNS_PRIME_BITS'd767637189, `RNS_PRIME_BITS'd847592127, `RNS_PRIME_BITS'd1721664702, `RNS_PRIME_BITS'd989079718, `RNS_PRIME_BITS'd1516681323},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd714854665, `RNS_PRIME_BITS'd133209267, `RNS_PRIME_BITS'd1030890025, `RNS_PRIME_BITS'd1797319518, `RNS_PRIME_BITS'd920238926, `RNS_PRIME_BITS'd468507401, `RNS_PRIME_BITS'd1476676690, `RNS_PRIME_BITS'd634956408, `RNS_PRIME_BITS'd1792572560, `RNS_PRIME_BITS'd61990415},
			'{`RNS_PRIME_BITS'd38, `RNS_PRIME_BITS'd1221081206, `RNS_PRIME_BITS'd563779542, `RNS_PRIME_BITS'd2030800400, `RNS_PRIME_BITS'd751293144, `RNS_PRIME_BITS'd229327497, `RNS_PRIME_BITS'd227263179, `RNS_PRIME_BITS'd1851316945, `RNS_PRIME_BITS'd732758559, `RNS_PRIME_BITS'd1593227780, `RNS_PRIME_BITS'd587733985},
			'{`RNS_PRIME_BITS'd191, `RNS_PRIME_BITS'd1807910007, `RNS_PRIME_BITS'd1619895485, `RNS_PRIME_BITS'd620061480, `RNS_PRIME_BITS'd768807831, `RNS_PRIME_BITS'd917985559, `RNS_PRIME_BITS'd1503055649, `RNS_PRIME_BITS'd719963627, `RNS_PRIME_BITS'd1472904887, `RNS_PRIME_BITS'd1581589716, `RNS_PRIME_BITS'd1439858118},
			'{`RNS_PRIME_BITS'd168, `RNS_PRIME_BITS'd1154482483, `RNS_PRIME_BITS'd1207323888, `RNS_PRIME_BITS'd1867975269, `RNS_PRIME_BITS'd1325265687, `RNS_PRIME_BITS'd600060113, `RNS_PRIME_BITS'd833046423, `RNS_PRIME_BITS'd41431813, `RNS_PRIME_BITS'd1659914147, `RNS_PRIME_BITS'd1016349382, `RNS_PRIME_BITS'd1508281587}
		},
		'{
			'{`RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd1955536273, `RNS_PRIME_BITS'd72199769, `RNS_PRIME_BITS'd543738865, `RNS_PRIME_BITS'd278149069, `RNS_PRIME_BITS'd112039133, `RNS_PRIME_BITS'd1423440261, `RNS_PRIME_BITS'd817119305, `RNS_PRIME_BITS'd96854077, `RNS_PRIME_BITS'd136144379, `RNS_PRIME_BITS'd290068202},
			'{`RNS_PRIME_BITS'd140, `RNS_PRIME_BITS'd1163932468, `RNS_PRIME_BITS'd1312115868, `RNS_PRIME_BITS'd1671692522, `RNS_PRIME_BITS'd413219362, `RNS_PRIME_BITS'd1713380497, `RNS_PRIME_BITS'd1617337393, `RNS_PRIME_BITS'd1825393305, `RNS_PRIME_BITS'd543164807, `RNS_PRIME_BITS'd174174202, `RNS_PRIME_BITS'd1617225077},
			'{`RNS_PRIME_BITS'd110, `RNS_PRIME_BITS'd1242824150, `RNS_PRIME_BITS'd1772024162, `RNS_PRIME_BITS'd1544376461, `RNS_PRIME_BITS'd1262406836, `RNS_PRIME_BITS'd847713700, `RNS_PRIME_BITS'd1793982018, `RNS_PRIME_BITS'd1650481697, `RNS_PRIME_BITS'd1529911082, `RNS_PRIME_BITS'd649737925, `RNS_PRIME_BITS'd1318527987},
			'{`RNS_PRIME_BITS'd107, `RNS_PRIME_BITS'd310553732, `RNS_PRIME_BITS'd965135146, `RNS_PRIME_BITS'd929301015, `RNS_PRIME_BITS'd277100629, `RNS_PRIME_BITS'd1079084040, `RNS_PRIME_BITS'd142532914, `RNS_PRIME_BITS'd599029720, `RNS_PRIME_BITS'd189404279, `RNS_PRIME_BITS'd1361295591, `RNS_PRIME_BITS'd1273942648},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1717285756, `RNS_PRIME_BITS'd2120818968, `RNS_PRIME_BITS'd413689768, `RNS_PRIME_BITS'd356200188, `RNS_PRIME_BITS'd965145043, `RNS_PRIME_BITS'd947752723, `RNS_PRIME_BITS'd1112660210, `RNS_PRIME_BITS'd693476553, `RNS_PRIME_BITS'd1461887076, `RNS_PRIME_BITS'd1014121477},
			'{`RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd1085810113, `RNS_PRIME_BITS'd2024319299, `RNS_PRIME_BITS'd1368882161, `RNS_PRIME_BITS'd903003222, `RNS_PRIME_BITS'd613533095, `RNS_PRIME_BITS'd363874595, `RNS_PRIME_BITS'd499314849, `RNS_PRIME_BITS'd1268597761, `RNS_PRIME_BITS'd1731796390, `RNS_PRIME_BITS'd260830956},
			'{`RNS_PRIME_BITS'd182, `RNS_PRIME_BITS'd589867125, `RNS_PRIME_BITS'd1767925930, `RNS_PRIME_BITS'd1491541114, `RNS_PRIME_BITS'd293741262, `RNS_PRIME_BITS'd1860795667, `RNS_PRIME_BITS'd2110253304, `RNS_PRIME_BITS'd512652926, `RNS_PRIME_BITS'd322295516, `RNS_PRIME_BITS'd881651729, `RNS_PRIME_BITS'd297248988},
			'{`RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd2047205371, `RNS_PRIME_BITS'd1369727446, `RNS_PRIME_BITS'd961432504, `RNS_PRIME_BITS'd607332966, `RNS_PRIME_BITS'd1082750757, `RNS_PRIME_BITS'd97009736, `RNS_PRIME_BITS'd856767739, `RNS_PRIME_BITS'd145039768, `RNS_PRIME_BITS'd11811546, `RNS_PRIME_BITS'd1138992481},
			'{`RNS_PRIME_BITS'd156, `RNS_PRIME_BITS'd283952402, `RNS_PRIME_BITS'd13218497, `RNS_PRIME_BITS'd1193417700, `RNS_PRIME_BITS'd232555216, `RNS_PRIME_BITS'd1788305925, `RNS_PRIME_BITS'd1733493902, `RNS_PRIME_BITS'd797373016, `RNS_PRIME_BITS'd224794926, `RNS_PRIME_BITS'd1326450227, `RNS_PRIME_BITS'd541377545},
			'{`RNS_PRIME_BITS'd19, `RNS_PRIME_BITS'd311191428, `RNS_PRIME_BITS'd1766396182, `RNS_PRIME_BITS'd106710594, `RNS_PRIME_BITS'd1383647258, `RNS_PRIME_BITS'd243603280, `RNS_PRIME_BITS'd361527932, `RNS_PRIME_BITS'd2092979402, `RNS_PRIME_BITS'd1708691588, `RNS_PRIME_BITS'd988480545, `RNS_PRIME_BITS'd722666355},
			'{`RNS_PRIME_BITS'd112, `RNS_PRIME_BITS'd1995201589, `RNS_PRIME_BITS'd1941322107, `RNS_PRIME_BITS'd2140276072, `RNS_PRIME_BITS'd1197697332, `RNS_PRIME_BITS'd388756108, `RNS_PRIME_BITS'd330686931, `RNS_PRIME_BITS'd73377547, `RNS_PRIME_BITS'd152624853, `RNS_PRIME_BITS'd491685070, `RNS_PRIME_BITS'd1554332703},
			'{`RNS_PRIME_BITS'd233, `RNS_PRIME_BITS'd670233579, `RNS_PRIME_BITS'd169768881, `RNS_PRIME_BITS'd2111380823, `RNS_PRIME_BITS'd472200319, `RNS_PRIME_BITS'd1739323043, `RNS_PRIME_BITS'd320644118, `RNS_PRIME_BITS'd1492857345, `RNS_PRIME_BITS'd821418206, `RNS_PRIME_BITS'd1983375056, `RNS_PRIME_BITS'd2117709478},
			'{`RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd1632926435, `RNS_PRIME_BITS'd417111103, `RNS_PRIME_BITS'd1298778681, `RNS_PRIME_BITS'd736680021, `RNS_PRIME_BITS'd1944265860, `RNS_PRIME_BITS'd1224087572, `RNS_PRIME_BITS'd1074246437, `RNS_PRIME_BITS'd1900343197, `RNS_PRIME_BITS'd1626925347, `RNS_PRIME_BITS'd1167086974},
			'{`RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd886535920, `RNS_PRIME_BITS'd1761969137, `RNS_PRIME_BITS'd60961537, `RNS_PRIME_BITS'd1971834382, `RNS_PRIME_BITS'd675730619, `RNS_PRIME_BITS'd1550400038, `RNS_PRIME_BITS'd1858681526, `RNS_PRIME_BITS'd315384538, `RNS_PRIME_BITS'd670869826, `RNS_PRIME_BITS'd484129533},
			'{`RNS_PRIME_BITS'd39, `RNS_PRIME_BITS'd1987160438, `RNS_PRIME_BITS'd697494481, `RNS_PRIME_BITS'd1740554836, `RNS_PRIME_BITS'd891344131, `RNS_PRIME_BITS'd1145005528, `RNS_PRIME_BITS'd1167416481, `RNS_PRIME_BITS'd1867470027, `RNS_PRIME_BITS'd1404495068, `RNS_PRIME_BITS'd204985604, `RNS_PRIME_BITS'd683670824},
			'{`RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd1281635686, `RNS_PRIME_BITS'd1934026553, `RNS_PRIME_BITS'd288726467, `RNS_PRIME_BITS'd527843471, `RNS_PRIME_BITS'd1094613239, `RNS_PRIME_BITS'd1740159566, `RNS_PRIME_BITS'd556004217, `RNS_PRIME_BITS'd670174587, `RNS_PRIME_BITS'd681185455, `RNS_PRIME_BITS'd408016772},
			'{`RNS_PRIME_BITS'd151, `RNS_PRIME_BITS'd2084195698, `RNS_PRIME_BITS'd1513483558, `RNS_PRIME_BITS'd735420047, `RNS_PRIME_BITS'd1352501917, `RNS_PRIME_BITS'd1700541820, `RNS_PRIME_BITS'd118030553, `RNS_PRIME_BITS'd351965771, `RNS_PRIME_BITS'd1516490344, `RNS_PRIME_BITS'd1342444826, `RNS_PRIME_BITS'd735768927},
			'{`RNS_PRIME_BITS'd53, `RNS_PRIME_BITS'd310971118, `RNS_PRIME_BITS'd756476479, `RNS_PRIME_BITS'd1855667466, `RNS_PRIME_BITS'd539151301, `RNS_PRIME_BITS'd1416767556, `RNS_PRIME_BITS'd1163136607, `RNS_PRIME_BITS'd1839074881, `RNS_PRIME_BITS'd1061101669, `RNS_PRIME_BITS'd1597184826, `RNS_PRIME_BITS'd649429200},
			'{`RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd1006915154, `RNS_PRIME_BITS'd361249612, `RNS_PRIME_BITS'd809079665, `RNS_PRIME_BITS'd2002997204, `RNS_PRIME_BITS'd1853846756, `RNS_PRIME_BITS'd943537268, `RNS_PRIME_BITS'd356909091, `RNS_PRIME_BITS'd1571400458, `RNS_PRIME_BITS'd1354755402, `RNS_PRIME_BITS'd49759249},
			'{`RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd1546481497, `RNS_PRIME_BITS'd302559892, `RNS_PRIME_BITS'd1410432228, `RNS_PRIME_BITS'd1506127415, `RNS_PRIME_BITS'd1583908025, `RNS_PRIME_BITS'd1988951365, `RNS_PRIME_BITS'd1512116038, `RNS_PRIME_BITS'd927402907, `RNS_PRIME_BITS'd1775440897, `RNS_PRIME_BITS'd979212807},
			'{`RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd1415549978, `RNS_PRIME_BITS'd683785885, `RNS_PRIME_BITS'd2116635297, `RNS_PRIME_BITS'd1092329007, `RNS_PRIME_BITS'd1914804675, `RNS_PRIME_BITS'd725064156, `RNS_PRIME_BITS'd1908636859, `RNS_PRIME_BITS'd1635625950, `RNS_PRIME_BITS'd1827207067, `RNS_PRIME_BITS'd1066563667},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1292288523, `RNS_PRIME_BITS'd35657733, `RNS_PRIME_BITS'd281361022, `RNS_PRIME_BITS'd726011793, `RNS_PRIME_BITS'd1075155106, `RNS_PRIME_BITS'd584885645, `RNS_PRIME_BITS'd1988349837, `RNS_PRIME_BITS'd915945215, `RNS_PRIME_BITS'd60981741, `RNS_PRIME_BITS'd2076342731},
			'{`RNS_PRIME_BITS'd119, `RNS_PRIME_BITS'd1615723254, `RNS_PRIME_BITS'd1106231901, `RNS_PRIME_BITS'd406084317, `RNS_PRIME_BITS'd501351162, `RNS_PRIME_BITS'd629266611, `RNS_PRIME_BITS'd907020161, `RNS_PRIME_BITS'd1228814670, `RNS_PRIME_BITS'd1287045125, `RNS_PRIME_BITS'd1001099801, `RNS_PRIME_BITS'd1373997896},
			'{`RNS_PRIME_BITS'd213, `RNS_PRIME_BITS'd491135873, `RNS_PRIME_BITS'd1918606366, `RNS_PRIME_BITS'd244259390, `RNS_PRIME_BITS'd1519001639, `RNS_PRIME_BITS'd1762335828, `RNS_PRIME_BITS'd360360711, `RNS_PRIME_BITS'd1779327718, `RNS_PRIME_BITS'd950511526, `RNS_PRIME_BITS'd1289223952, `RNS_PRIME_BITS'd2061738439},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd2115206369, `RNS_PRIME_BITS'd832381212, `RNS_PRIME_BITS'd1258227420, `RNS_PRIME_BITS'd240051297, `RNS_PRIME_BITS'd1176235920, `RNS_PRIME_BITS'd1368868271, `RNS_PRIME_BITS'd2055487246, `RNS_PRIME_BITS'd87511821, `RNS_PRIME_BITS'd1598504741, `RNS_PRIME_BITS'd1079748956},
			'{`RNS_PRIME_BITS'd7, `RNS_PRIME_BITS'd2020287580, `RNS_PRIME_BITS'd1067618791, `RNS_PRIME_BITS'd113597757, `RNS_PRIME_BITS'd1393196806, `RNS_PRIME_BITS'd196447480, `RNS_PRIME_BITS'd327922108, `RNS_PRIME_BITS'd1759803643, `RNS_PRIME_BITS'd1931942087, `RNS_PRIME_BITS'd13870182, `RNS_PRIME_BITS'd959307838},
			'{`RNS_PRIME_BITS'd104, `RNS_PRIME_BITS'd1914429170, `RNS_PRIME_BITS'd223667310, `RNS_PRIME_BITS'd948402256, `RNS_PRIME_BITS'd1915142970, `RNS_PRIME_BITS'd150135089, `RNS_PRIME_BITS'd490224957, `RNS_PRIME_BITS'd1313831840, `RNS_PRIME_BITS'd484922740, `RNS_PRIME_BITS'd1087821508, `RNS_PRIME_BITS'd754973320},
			'{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd2102216063, `RNS_PRIME_BITS'd1837188824, `RNS_PRIME_BITS'd1669094389, `RNS_PRIME_BITS'd1118969516, `RNS_PRIME_BITS'd1745612743, `RNS_PRIME_BITS'd1856426117, `RNS_PRIME_BITS'd1662497348, `RNS_PRIME_BITS'd2059035398, `RNS_PRIME_BITS'd1840250640, `RNS_PRIME_BITS'd1845798413},
			'{`RNS_PRIME_BITS'd63, `RNS_PRIME_BITS'd2004737626, `RNS_PRIME_BITS'd2108414541, `RNS_PRIME_BITS'd369794248, `RNS_PRIME_BITS'd878244132, `RNS_PRIME_BITS'd626065828, `RNS_PRIME_BITS'd2063810886, `RNS_PRIME_BITS'd2007244949, `RNS_PRIME_BITS'd2008923671, `RNS_PRIME_BITS'd1242808099, `RNS_PRIME_BITS'd513565533},
			'{`RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd1137118902, `RNS_PRIME_BITS'd872008029, `RNS_PRIME_BITS'd191416066, `RNS_PRIME_BITS'd62240418, `RNS_PRIME_BITS'd413727601, `RNS_PRIME_BITS'd1248446497, `RNS_PRIME_BITS'd460803719, `RNS_PRIME_BITS'd1409848599, `RNS_PRIME_BITS'd108429392, `RNS_PRIME_BITS'd1565502727},
			'{`RNS_PRIME_BITS'd41, `RNS_PRIME_BITS'd486757631, `RNS_PRIME_BITS'd428774361, `RNS_PRIME_BITS'd1444831977, `RNS_PRIME_BITS'd935428476, `RNS_PRIME_BITS'd719923345, `RNS_PRIME_BITS'd941058696, `RNS_PRIME_BITS'd689636971, `RNS_PRIME_BITS'd229607187, `RNS_PRIME_BITS'd377792345, `RNS_PRIME_BITS'd145157527},
			'{`RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd382599106, `RNS_PRIME_BITS'd1942241138, `RNS_PRIME_BITS'd1511641449, `RNS_PRIME_BITS'd101951284, `RNS_PRIME_BITS'd755762491, `RNS_PRIME_BITS'd1393396211, `RNS_PRIME_BITS'd987108858, `RNS_PRIME_BITS'd850982833, `RNS_PRIME_BITS'd1067316770, `RNS_PRIME_BITS'd1808764233},
			'{`RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd1532552119, `RNS_PRIME_BITS'd835413317, `RNS_PRIME_BITS'd62466030, `RNS_PRIME_BITS'd1471861893, `RNS_PRIME_BITS'd141765467, `RNS_PRIME_BITS'd1959625611, `RNS_PRIME_BITS'd1079664426, `RNS_PRIME_BITS'd803942275, `RNS_PRIME_BITS'd2054128965, `RNS_PRIME_BITS'd1874294153},
			'{`RNS_PRIME_BITS'd48, `RNS_PRIME_BITS'd737416758, `RNS_PRIME_BITS'd1430247446, `RNS_PRIME_BITS'd748173331, `RNS_PRIME_BITS'd1074972251, `RNS_PRIME_BITS'd754076283, `RNS_PRIME_BITS'd348148591, `RNS_PRIME_BITS'd454414574, `RNS_PRIME_BITS'd1040205047, `RNS_PRIME_BITS'd809995724, `RNS_PRIME_BITS'd1309216869},
			'{`RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd1064729691, `RNS_PRIME_BITS'd277424839, `RNS_PRIME_BITS'd1187108361, `RNS_PRIME_BITS'd1892974459, `RNS_PRIME_BITS'd794803551, `RNS_PRIME_BITS'd2056766307, `RNS_PRIME_BITS'd959428892, `RNS_PRIME_BITS'd839775371, `RNS_PRIME_BITS'd1353166206, `RNS_PRIME_BITS'd48585900},
			'{`RNS_PRIME_BITS'd221, `RNS_PRIME_BITS'd1969409989, `RNS_PRIME_BITS'd502890567, `RNS_PRIME_BITS'd1617498340, `RNS_PRIME_BITS'd268326264, `RNS_PRIME_BITS'd739247882, `RNS_PRIME_BITS'd1976574944, `RNS_PRIME_BITS'd828259338, `RNS_PRIME_BITS'd1873743871, `RNS_PRIME_BITS'd1046172520, `RNS_PRIME_BITS'd916356759},
			'{`RNS_PRIME_BITS'd160, `RNS_PRIME_BITS'd1302474013, `RNS_PRIME_BITS'd2122105034, `RNS_PRIME_BITS'd767262510, `RNS_PRIME_BITS'd325521869, `RNS_PRIME_BITS'd185538554, `RNS_PRIME_BITS'd969860449, `RNS_PRIME_BITS'd315169130, `RNS_PRIME_BITS'd1952047749, `RNS_PRIME_BITS'd774280044, `RNS_PRIME_BITS'd930177179},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd119967844, `RNS_PRIME_BITS'd2143443333, `RNS_PRIME_BITS'd1465877926, `RNS_PRIME_BITS'd89512082, `RNS_PRIME_BITS'd241598987, `RNS_PRIME_BITS'd1082821552, `RNS_PRIME_BITS'd2025769303, `RNS_PRIME_BITS'd1971415449, `RNS_PRIME_BITS'd1507042086, `RNS_PRIME_BITS'd692338999},
			'{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd1808660323, `RNS_PRIME_BITS'd1890233008, `RNS_PRIME_BITS'd908191028, `RNS_PRIME_BITS'd858820278, `RNS_PRIME_BITS'd1527453734, `RNS_PRIME_BITS'd864766317, `RNS_PRIME_BITS'd1419049821, `RNS_PRIME_BITS'd1096040475, `RNS_PRIME_BITS'd492638349, `RNS_PRIME_BITS'd1127659372},
			'{`RNS_PRIME_BITS'd166, `RNS_PRIME_BITS'd214998419, `RNS_PRIME_BITS'd232816601, `RNS_PRIME_BITS'd1980306491, `RNS_PRIME_BITS'd424502640, `RNS_PRIME_BITS'd398490968, `RNS_PRIME_BITS'd36859219, `RNS_PRIME_BITS'd546651679, `RNS_PRIME_BITS'd489724868, `RNS_PRIME_BITS'd1519270358, `RNS_PRIME_BITS'd1009311657},
			'{`RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd2106270946, `RNS_PRIME_BITS'd1641208426, `RNS_PRIME_BITS'd277748957, `RNS_PRIME_BITS'd1411464231, `RNS_PRIME_BITS'd2116615443, `RNS_PRIME_BITS'd2062845646, `RNS_PRIME_BITS'd11316339, `RNS_PRIME_BITS'd1761931607, `RNS_PRIME_BITS'd1652274179, `RNS_PRIME_BITS'd1905135075},
			'{`RNS_PRIME_BITS'd10, `RNS_PRIME_BITS'd1483702020, `RNS_PRIME_BITS'd528311709, `RNS_PRIME_BITS'd1962963232, `RNS_PRIME_BITS'd966507989, `RNS_PRIME_BITS'd2134090138, `RNS_PRIME_BITS'd1037191895, `RNS_PRIME_BITS'd373746857, `RNS_PRIME_BITS'd1857699132, `RNS_PRIME_BITS'd1536659203, `RNS_PRIME_BITS'd92773432},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd693731814, `RNS_PRIME_BITS'd111629882, `RNS_PRIME_BITS'd1714436560, `RNS_PRIME_BITS'd1464101822, `RNS_PRIME_BITS'd1597965284, `RNS_PRIME_BITS'd1448580154, `RNS_PRIME_BITS'd1403549376, `RNS_PRIME_BITS'd1403949919, `RNS_PRIME_BITS'd1189412705, `RNS_PRIME_BITS'd1853813266},
			'{`RNS_PRIME_BITS'd214, `RNS_PRIME_BITS'd556136742, `RNS_PRIME_BITS'd936666090, `RNS_PRIME_BITS'd1401073343, `RNS_PRIME_BITS'd1438355215, `RNS_PRIME_BITS'd554106083, `RNS_PRIME_BITS'd63923294, `RNS_PRIME_BITS'd1768110488, `RNS_PRIME_BITS'd583359313, `RNS_PRIME_BITS'd853101852, `RNS_PRIME_BITS'd1125956773},
			'{`RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd1629132477, `RNS_PRIME_BITS'd1490326907, `RNS_PRIME_BITS'd71237407, `RNS_PRIME_BITS'd2122676209, `RNS_PRIME_BITS'd1196265291, `RNS_PRIME_BITS'd673765066, `RNS_PRIME_BITS'd1560991675, `RNS_PRIME_BITS'd486425493, `RNS_PRIME_BITS'd1098046388, `RNS_PRIME_BITS'd1588331160},
			'{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd159875036, `RNS_PRIME_BITS'd949410008, `RNS_PRIME_BITS'd1223223189, `RNS_PRIME_BITS'd1217243037, `RNS_PRIME_BITS'd2134785112, `RNS_PRIME_BITS'd339782542, `RNS_PRIME_BITS'd1753210772, `RNS_PRIME_BITS'd378401668, `RNS_PRIME_BITS'd1033418253, `RNS_PRIME_BITS'd25930037},
			'{`RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd148909854, `RNS_PRIME_BITS'd69349500, `RNS_PRIME_BITS'd1103780858, `RNS_PRIME_BITS'd829179584, `RNS_PRIME_BITS'd1560313955, `RNS_PRIME_BITS'd1685953918, `RNS_PRIME_BITS'd1957316237, `RNS_PRIME_BITS'd1651498874, `RNS_PRIME_BITS'd929139619, `RNS_PRIME_BITS'd336392472},
			'{`RNS_PRIME_BITS'd106, `RNS_PRIME_BITS'd1418329607, `RNS_PRIME_BITS'd2146952119, `RNS_PRIME_BITS'd1421992412, `RNS_PRIME_BITS'd732950140, `RNS_PRIME_BITS'd1424849677, `RNS_PRIME_BITS'd1602557241, `RNS_PRIME_BITS'd72626322, `RNS_PRIME_BITS'd1119580274, `RNS_PRIME_BITS'd330998865, `RNS_PRIME_BITS'd1671958619},
			'{`RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd522561120, `RNS_PRIME_BITS'd665745394, `RNS_PRIME_BITS'd278258742, `RNS_PRIME_BITS'd736709169, `RNS_PRIME_BITS'd1155273371, `RNS_PRIME_BITS'd980637863, `RNS_PRIME_BITS'd2030774306, `RNS_PRIME_BITS'd4198333, `RNS_PRIME_BITS'd950911550, `RNS_PRIME_BITS'd421474428},
			'{`RNS_PRIME_BITS'd78, `RNS_PRIME_BITS'd306753226, `RNS_PRIME_BITS'd438693194, `RNS_PRIME_BITS'd375058046, `RNS_PRIME_BITS'd1849117976, `RNS_PRIME_BITS'd1382746700, `RNS_PRIME_BITS'd587982605, `RNS_PRIME_BITS'd695777053, `RNS_PRIME_BITS'd1405502169, `RNS_PRIME_BITS'd120180029, `RNS_PRIME_BITS'd271779404},
			'{`RNS_PRIME_BITS'd181, `RNS_PRIME_BITS'd649796929, `RNS_PRIME_BITS'd863617473, `RNS_PRIME_BITS'd23649474, `RNS_PRIME_BITS'd1104446652, `RNS_PRIME_BITS'd1017117469, `RNS_PRIME_BITS'd593514738, `RNS_PRIME_BITS'd1070307677, `RNS_PRIME_BITS'd409010570, `RNS_PRIME_BITS'd825464853, `RNS_PRIME_BITS'd1037680112},
			'{`RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd195647729, `RNS_PRIME_BITS'd1063252121, `RNS_PRIME_BITS'd1538741575, `RNS_PRIME_BITS'd2123704085, `RNS_PRIME_BITS'd161471826, `RNS_PRIME_BITS'd299831853, `RNS_PRIME_BITS'd91222297, `RNS_PRIME_BITS'd1861375948, `RNS_PRIME_BITS'd1765379990, `RNS_PRIME_BITS'd744565894},
			'{`RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd981115086, `RNS_PRIME_BITS'd1188660595, `RNS_PRIME_BITS'd332658162, `RNS_PRIME_BITS'd1047116775, `RNS_PRIME_BITS'd86592155, `RNS_PRIME_BITS'd1301046809, `RNS_PRIME_BITS'd969677079, `RNS_PRIME_BITS'd992504658, `RNS_PRIME_BITS'd1679087270, `RNS_PRIME_BITS'd931158969},
			'{`RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd367209162, `RNS_PRIME_BITS'd303848766, `RNS_PRIME_BITS'd1211880725, `RNS_PRIME_BITS'd1633199764, `RNS_PRIME_BITS'd755803528, `RNS_PRIME_BITS'd157436782, `RNS_PRIME_BITS'd546282529, `RNS_PRIME_BITS'd1608589642, `RNS_PRIME_BITS'd1546861089, `RNS_PRIME_BITS'd1741944937},
			'{`RNS_PRIME_BITS'd96, `RNS_PRIME_BITS'd393994442, `RNS_PRIME_BITS'd1893446090, `RNS_PRIME_BITS'd1168901681, `RNS_PRIME_BITS'd1329060816, `RNS_PRIME_BITS'd1079743521, `RNS_PRIME_BITS'd1377889218, `RNS_PRIME_BITS'd583181574, `RNS_PRIME_BITS'd1182907980, `RNS_PRIME_BITS'd460196244, `RNS_PRIME_BITS'd1888190241},
			'{`RNS_PRIME_BITS'd194, `RNS_PRIME_BITS'd169104737, `RNS_PRIME_BITS'd368323366, `RNS_PRIME_BITS'd1032409385, `RNS_PRIME_BITS'd479517844, `RNS_PRIME_BITS'd708821118, `RNS_PRIME_BITS'd911576691, `RNS_PRIME_BITS'd682948336, `RNS_PRIME_BITS'd2114988917, `RNS_PRIME_BITS'd423859014, `RNS_PRIME_BITS'd1931554656},
			'{`RNS_PRIME_BITS'd165, `RNS_PRIME_BITS'd1450489498, `RNS_PRIME_BITS'd1583408245, `RNS_PRIME_BITS'd407370474, `RNS_PRIME_BITS'd1463908530, `RNS_PRIME_BITS'd986483440, `RNS_PRIME_BITS'd1052436246, `RNS_PRIME_BITS'd510606176, `RNS_PRIME_BITS'd2014458801, `RNS_PRIME_BITS'd1266526573, `RNS_PRIME_BITS'd417574515},
			'{`RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd1797127746, `RNS_PRIME_BITS'd1728314843, `RNS_PRIME_BITS'd141522374, `RNS_PRIME_BITS'd265458872, `RNS_PRIME_BITS'd2016725951, `RNS_PRIME_BITS'd441876223, `RNS_PRIME_BITS'd651437286, `RNS_PRIME_BITS'd1479640758, `RNS_PRIME_BITS'd90398282, `RNS_PRIME_BITS'd2129364097},
			'{`RNS_PRIME_BITS'd103, `RNS_PRIME_BITS'd435909378, `RNS_PRIME_BITS'd1159301959, `RNS_PRIME_BITS'd1402648299, `RNS_PRIME_BITS'd1214699232, `RNS_PRIME_BITS'd603643622, `RNS_PRIME_BITS'd574971132, `RNS_PRIME_BITS'd102669563, `RNS_PRIME_BITS'd1070168481, `RNS_PRIME_BITS'd1408643251, `RNS_PRIME_BITS'd2121821680},
			'{`RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd883857597, `RNS_PRIME_BITS'd221607576, `RNS_PRIME_BITS'd1193421194, `RNS_PRIME_BITS'd1796680906, `RNS_PRIME_BITS'd777854019, `RNS_PRIME_BITS'd2118245076, `RNS_PRIME_BITS'd711686997, `RNS_PRIME_BITS'd1187624587, `RNS_PRIME_BITS'd976328176, `RNS_PRIME_BITS'd777946846},
			'{`RNS_PRIME_BITS'd183, `RNS_PRIME_BITS'd1907927343, `RNS_PRIME_BITS'd1428177263, `RNS_PRIME_BITS'd1915120244, `RNS_PRIME_BITS'd189443874, `RNS_PRIME_BITS'd668765619, `RNS_PRIME_BITS'd1887426247, `RNS_PRIME_BITS'd436714259, `RNS_PRIME_BITS'd1206207826, `RNS_PRIME_BITS'd150495050, `RNS_PRIME_BITS'd1473065914},
			'{`RNS_PRIME_BITS'd54, `RNS_PRIME_BITS'd62201952, `RNS_PRIME_BITS'd1586795134, `RNS_PRIME_BITS'd413919165, `RNS_PRIME_BITS'd1804883783, `RNS_PRIME_BITS'd199655685, `RNS_PRIME_BITS'd1232564150, `RNS_PRIME_BITS'd1009449661, `RNS_PRIME_BITS'd141185226, `RNS_PRIME_BITS'd981792410, `RNS_PRIME_BITS'd644083540},
			'{`RNS_PRIME_BITS'd82, `RNS_PRIME_BITS'd1282705513, `RNS_PRIME_BITS'd831740344, `RNS_PRIME_BITS'd1680158077, `RNS_PRIME_BITS'd1862197948, `RNS_PRIME_BITS'd1072876092, `RNS_PRIME_BITS'd1419289202, `RNS_PRIME_BITS'd2070584480, `RNS_PRIME_BITS'd1678758297, `RNS_PRIME_BITS'd218302214, `RNS_PRIME_BITS'd536262211},
			'{`RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd322917985, `RNS_PRIME_BITS'd1096008895, `RNS_PRIME_BITS'd1082599150, `RNS_PRIME_BITS'd299744371, `RNS_PRIME_BITS'd1021539026, `RNS_PRIME_BITS'd2032943338, `RNS_PRIME_BITS'd445874010, `RNS_PRIME_BITS'd477550301, `RNS_PRIME_BITS'd1562517956, `RNS_PRIME_BITS'd1395797683}
		}
	}
};


// ---------------------------
// Operation/Control Types & misc
// ---------------------------

// how many polynomials can the register file store
`define REG_NPOLY 12

// If you ever want to explicitly tag A vs B in code:
typedef enum logic [0:0] {
  POLY_A = 1'b0,
  POLY_B = 1'b1
} poly_sel_e;

typedef enum logic [2:0] {
    NO_OP,
    OP_CT_CT_ADD,
    OP_CT_PT_ADD,
    OP_CT_PT_MUL,
    OP_CT_CT_MUL
} op_e;

typedef struct packed {
  op_e                          mode;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_b;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_b;
  logic [$clog2(`REG_NPOLY)-1:0]      out_a;
  logic [$clog2(`REG_NPOLY)-1:0]      out_b;
} operation;

// program counter (aka current state) is 5 bits = up to 32 states
`define PROGRAM_COUNTER_BITS 7
typedef logic [`PROGRAM_COUNTER_BITS-1:0] pc_state_type; 

`endif
