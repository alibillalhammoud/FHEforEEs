`ifndef TYPES_SVH
`define TYPES_SVH

// ---------------------------
// Basic data types
// ---------------------------



// NTT
`define BASE      32'd2
// Width of each RNS residue (one small prime)
`define RNS_PRIME_BITS 32
// RNS residues
typedef logic [`RNS_PRIME_BITS-1:0] rns_residue_t; 
typedef logic [(2*`RNS_PRIME_BITS)-1:0] wide_rns_residue_t;
// Vector / slot params
`define N_SLOTS   64
// moduli and RNS bases
`define t_MODULUS 257

`define q_BASIS_LEN 11
//`define q_MODULUS = 536092687689737712660299305370020840707037344303743567681198293980556215074372863278673727266177
parameter rns_residue_t q_BASIS [`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353};
//`define B_MODULUS = 2086045702160390514072457421164142647843268814746900546792219301529141418454085790414389880321
`define B_BASIS_LEN 10
parameter rns_residue_t B_BASIS [`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337};
//`define Ba_MODULUS = 2147503489
`define Ba_BASIS_LEN 1
parameter rns_residue_t Ba_BASIS [`Ba_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147503489};
`define qBBa_BASIS_LEN 22
//`define qBBa_MODULUS = 2401582888476023779443294070753805757615044045174800139284098902756577490274881128570727198734820745298450301532339857214864378319647024214690248526201090429246246041638715397173165827069546764128513
parameter rns_residue_t qBBa_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd257, `RNS_PRIME_BITS'd2147483777, `RNS_PRIME_BITS'd2147484161, `RNS_PRIME_BITS'd2147484929, `RNS_PRIME_BITS'd2147485057, `RNS_PRIME_BITS'd2147486849, `RNS_PRIME_BITS'd2147488001, `RNS_PRIME_BITS'd2147489537, `RNS_PRIME_BITS'd2147490689, `RNS_PRIME_BITS'd2147491201, `RNS_PRIME_BITS'd2147492353, `RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147503489};
parameter rns_residue_t w_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd1684230034, `RNS_PRIME_BITS'd413528229, `RNS_PRIME_BITS'd835068854, `RNS_PRIME_BITS'd698897645, `RNS_PRIME_BITS'd266488565, `RNS_PRIME_BITS'd1915797300, `RNS_PRIME_BITS'd634442553, `RNS_PRIME_BITS'd207695132, `RNS_PRIME_BITS'd21725588, `RNS_PRIME_BITS'd209219715, `RNS_PRIME_BITS'd1654849230, `RNS_PRIME_BITS'd318222520, `RNS_PRIME_BITS'd458644985, `RNS_PRIME_BITS'd1659477478, `RNS_PRIME_BITS'd221897449, `RNS_PRIME_BITS'd1817702166, `RNS_PRIME_BITS'd1453892451, `RNS_PRIME_BITS'd1033346514, `RNS_PRIME_BITS'd1445995283, `RNS_PRIME_BITS'd330138710, `RNS_PRIME_BITS'd545722081};
parameter rns_residue_t w_INV_BASIS [`qBBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd165, `RNS_PRIME_BITS'd465883484, `RNS_PRIME_BITS'd1309966555, `RNS_PRIME_BITS'd1089826325, `RNS_PRIME_BITS'd123767386, `RNS_PRIME_BITS'd1570352642, `RNS_PRIME_BITS'd374598187, `RNS_PRIME_BITS'd199676388, `RNS_PRIME_BITS'd1965833606, `RNS_PRIME_BITS'd1344902099, `RNS_PRIME_BITS'd1350503019, `RNS_PRIME_BITS'd1320961193, `RNS_PRIME_BITS'd1595145660, `RNS_PRIME_BITS'd673021473, `RNS_PRIME_BITS'd1565830187, `RNS_PRIME_BITS'd46526017, `RNS_PRIME_BITS'd1553448153, `RNS_PRIME_BITS'd1394618113, `RNS_PRIME_BITS'd1852124673, `RNS_PRIME_BITS'd1285194286, `RNS_PRIME_BITS'd438577756, `RNS_PRIME_BITS'd433881419};

`define BBa_BASIS_LEN 11
parameter rns_residue_t BBa_BASIS [`BBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd2147492609, `RNS_PRIME_BITS'd2147493889, `RNS_PRIME_BITS'd2147494273, `RNS_PRIME_BITS'd2147494529, `RNS_PRIME_BITS'd2147494913, `RNS_PRIME_BITS'd2147495681, `RNS_PRIME_BITS'd2147496193, `RNS_PRIME_BITS'd2147496961, `RNS_PRIME_BITS'd2147499521, `RNS_PRIME_BITS'd2147502337, `RNS_PRIME_BITS'd2147503489};

// RNS integers
typedef rns_residue_t rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef rns_residue_t rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef rns_residue_t rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
/*typedef rns_residue_t rns_coef_qBBa_BASIS_t [`q_BASIS_LEN + `B_BASIS_LEN + `Ba_BASIS_LEN];*/
// Polynomials
typedef rns_int_q_BASIS_t q_BASIS_poly [`N_SLOTS]; // 
typedef rns_int_B_BASIS_t B_BASIS_poly [`N_SLOTS]; //  
typedef rns_int_Ba_BASIS_t Ba_BASIS_poly [`N_SLOTS];
/*typedef rns_coef_qBBA_BASIS_t qBBa_BASIS_poly [`N_SLOTS];*/
// wide RNS integers (each residue is double the length for mult)
typedef wide_rns_residue_t wide_rns_int_q_BASIS_t [`q_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_B_BASIS_t [`B_BASIS_LEN];
typedef wide_rns_residue_t wide_rns_int_Ba_BASIS_t [`Ba_BASIS_LEN];
// wide Polynomials
typedef wide_rns_int_q_BASIS_t wide_q_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_B_BASIS_t wide_B_BASIS_poly [`N_SLOTS];
typedef wide_rns_int_Ba_BASIS_t wide_Ba_BASIS_poly [`N_SLOTS];

// ---------------------------
// precalculated values
// ---------------------------
// Example constant “twist” factors (all 1s for now)
parameter q_BASIS_poly twist_factor_q   = '{
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd9, `RNS_PRIME_BITS'd81, `RNS_PRIME_BITS'd215, `RNS_PRIME_BITS'd136, `RNS_PRIME_BITS'd196, `RNS_PRIME_BITS'd222, `RNS_PRIME_BITS'd199, `RNS_PRIME_BITS'd249, `RNS_PRIME_BITS'd185, `RNS_PRIME_BITS'd123, `RNS_PRIME_BITS'd79, `RNS_PRIME_BITS'd197, `RNS_PRIME_BITS'd231, `RNS_PRIME_BITS'd23, `RNS_PRIME_BITS'd207, `RNS_PRIME_BITS'd64, `RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd44, `RNS_PRIME_BITS'd139, `RNS_PRIME_BITS'd223, `RNS_PRIME_BITS'd208, `RNS_PRIME_BITS'd73, `RNS_PRIME_BITS'd143, `RNS_PRIME_BITS'd2, `RNS_PRIME_BITS'd18, `RNS_PRIME_BITS'd162, `RNS_PRIME_BITS'd173, `RNS_PRIME_BITS'd15, `RNS_PRIME_BITS'd135, `RNS_PRIME_BITS'd187, `RNS_PRIME_BITS'd141, `RNS_PRIME_BITS'd241, `RNS_PRIME_BITS'd113, `RNS_PRIME_BITS'd246, `RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd137, `RNS_PRIME_BITS'd205, `RNS_PRIME_BITS'd46, `RNS_PRIME_BITS'd157, `RNS_PRIME_BITS'd128, `RNS_PRIME_BITS'd124, `RNS_PRIME_BITS'd88, `RNS_PRIME_BITS'd21, `RNS_PRIME_BITS'd189, `RNS_PRIME_BITS'd159, `RNS_PRIME_BITS'd146, `RNS_PRIME_BITS'd29, `RNS_PRIME_BITS'd4, `RNS_PRIME_BITS'd36, `RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd57},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1454056114, `RNS_PRIME_BITS'd1684230034, `RNS_PRIME_BITS'd1874017521, `RNS_PRIME_BITS'd120548658, `RNS_PRIME_BITS'd340182173, `RNS_PRIME_BITS'd656530581, `RNS_PRIME_BITS'd1079385897, `RNS_PRIME_BITS'd1323801281, `RNS_PRIME_BITS'd1753733667, `RNS_PRIME_BITS'd109329595, `RNS_PRIME_BITS'd1102767568, `RNS_PRIME_BITS'd2066618854, `RNS_PRIME_BITS'd1323556320, `RNS_PRIME_BITS'd668212887, `RNS_PRIME_BITS'd1871724384, `RNS_PRIME_BITS'd1061363846, `RNS_PRIME_BITS'd248740266, `RNS_PRIME_BITS'd918758775, `RNS_PRIME_BITS'd1340620076, `RNS_PRIME_BITS'd1215568715, `RNS_PRIME_BITS'd16030913, `RNS_PRIME_BITS'd1583075798, `RNS_PRIME_BITS'd702020947, `RNS_PRIME_BITS'd426187835, `RNS_PRIME_BITS'd1577612670, `RNS_PRIME_BITS'd994527522, `RNS_PRIME_BITS'd994513885, `RNS_PRIME_BITS'd1896484085, `RNS_PRIME_BITS'd1390505442, `RNS_PRIME_BITS'd470517865, `RNS_PRIME_BITS'd1521041901, `RNS_PRIME_BITS'd1021707020, `RNS_PRIME_BITS'd774040236, `RNS_PRIME_BITS'd42370405, `RNS_PRIME_BITS'd1260414647, `RNS_PRIME_BITS'd2121222217, `RNS_PRIME_BITS'd1547276440, `RNS_PRIME_BITS'd1934841955, `RNS_PRIME_BITS'd883135528, `RNS_PRIME_BITS'd1146745373, `RNS_PRIME_BITS'd501271165, `RNS_PRIME_BITS'd788019979, `RNS_PRIME_BITS'd1009909057, `RNS_PRIME_BITS'd1963269275, `RNS_PRIME_BITS'd1270209618, `RNS_PRIME_BITS'd763626807, `RNS_PRIME_BITS'd480335015, `RNS_PRIME_BITS'd910119688, `RNS_PRIME_BITS'd1159872543, `RNS_PRIME_BITS'd1182896170, `RNS_PRIME_BITS'd350490837, `RNS_PRIME_BITS'd2086471810, `RNS_PRIME_BITS'd1074706051, `RNS_PRIME_BITS'd248908061, `RNS_PRIME_BITS'd42567327, `RNS_PRIME_BITS'd1605683, `RNS_PRIME_BITS'd231006354, `RNS_PRIME_BITS'd328404460, `RNS_PRIME_BITS'd184517896, `RNS_PRIME_BITS'd1628067296, `RNS_PRIME_BITS'd1495990324, `RNS_PRIME_BITS'd1681600293, `RNS_PRIME_BITS'd1180703254},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd2023476074, `RNS_PRIME_BITS'd413528229, `RNS_PRIME_BITS'd1276327416, `RNS_PRIME_BITS'd67511054, `RNS_PRIME_BITS'd951629099, `RNS_PRIME_BITS'd861227005, `RNS_PRIME_BITS'd576378926, `RNS_PRIME_BITS'd1485798473, `RNS_PRIME_BITS'd857515399, `RNS_PRIME_BITS'd1603393679, `RNS_PRIME_BITS'd1804390941, `RNS_PRIME_BITS'd1867409965, `RNS_PRIME_BITS'd2064658918, `RNS_PRIME_BITS'd1957088536, `RNS_PRIME_BITS'd1016906757, `RNS_PRIME_BITS'd2093569547, `RNS_PRIME_BITS'd1953159839, `RNS_PRIME_BITS'd74609970, `RNS_PRIME_BITS'd435782459, `RNS_PRIME_BITS'd764376413, `RNS_PRIME_BITS'd1073050120, `RNS_PRIME_BITS'd599521406, `RNS_PRIME_BITS'd1695639893, `RNS_PRIME_BITS'd1884145470, `RNS_PRIME_BITS'd1387757027, `RNS_PRIME_BITS'd837323404, `RNS_PRIME_BITS'd1449362922, `RNS_PRIME_BITS'd1456040658, `RNS_PRIME_BITS'd1703996997, `RNS_PRIME_BITS'd1343049929, `RNS_PRIME_BITS'd788800085, `RNS_PRIME_BITS'd434575099, `RNS_PRIME_BITS'd572591813, `RNS_PRIME_BITS'd813012214, `RNS_PRIME_BITS'd1319821704, `RNS_PRIME_BITS'd1458297369, `RNS_PRIME_BITS'd688415855, `RNS_PRIME_BITS'd34272266, `RNS_PRIME_BITS'd514568416, `RNS_PRIME_BITS'd108956348, `RNS_PRIME_BITS'd1695216211, `RNS_PRIME_BITS'd1530978778, `RNS_PRIME_BITS'd1563397195, `RNS_PRIME_BITS'd1871639102, `RNS_PRIME_BITS'd572522453, `RNS_PRIME_BITS'd1339861729, `RNS_PRIME_BITS'd800312580, `RNS_PRIME_BITS'd1128292512, `RNS_PRIME_BITS'd1784665556, `RNS_PRIME_BITS'd113138122, `RNS_PRIME_BITS'd228923992, `RNS_PRIME_BITS'd31790164, `RNS_PRIME_BITS'd183046999, `RNS_PRIME_BITS'd984227194, `RNS_PRIME_BITS'd1940067462, `RNS_PRIME_BITS'd397906100, `RNS_PRIME_BITS'd377036607, `RNS_PRIME_BITS'd1578585534, `RNS_PRIME_BITS'd1760756591, `RNS_PRIME_BITS'd445410876, `RNS_PRIME_BITS'd384884134, `RNS_PRIME_BITS'd837517606, `RNS_PRIME_BITS'd718232802},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1829761212, `RNS_PRIME_BITS'd835068854, `RNS_PRIME_BITS'd765723923, `RNS_PRIME_BITS'd346940440, `RNS_PRIME_BITS'd538002895, `RNS_PRIME_BITS'd1064440654, `RNS_PRIME_BITS'd1614098500, `RNS_PRIME_BITS'd469931230, `RNS_PRIME_BITS'd1345302327, `RNS_PRIME_BITS'd1699086710, `RNS_PRIME_BITS'd190235933, `RNS_PRIME_BITS'd973917268, `RNS_PRIME_BITS'd1573977587, `RNS_PRIME_BITS'd765942372, `RNS_PRIME_BITS'd631590787, `RNS_PRIME_BITS'd239311507, `RNS_PRIME_BITS'd793606413, `RNS_PRIME_BITS'd1368161792, `RNS_PRIME_BITS'd1256631702, `RNS_PRIME_BITS'd1968585711, `RNS_PRIME_BITS'd56850842, `RNS_PRIME_BITS'd2122922145, `RNS_PRIME_BITS'd1904384299, `RNS_PRIME_BITS'd514016804, `RNS_PRIME_BITS'd1634409210, `RNS_PRIME_BITS'd552952089, `RNS_PRIME_BITS'd257231880, `RNS_PRIME_BITS'd998069335, `RNS_PRIME_BITS'd132272763, `RNS_PRIME_BITS'd242912769, `RNS_PRIME_BITS'd185065907, `RNS_PRIME_BITS'd1712127733, `RNS_PRIME_BITS'd1210603202, `RNS_PRIME_BITS'd1479849359, `RNS_PRIME_BITS'd618256455, `RNS_PRIME_BITS'd336159836, `RNS_PRIME_BITS'd618238460, `RNS_PRIME_BITS'd1169566253, `RNS_PRIME_BITS'd1653743872, `RNS_PRIME_BITS'd230876332, `RNS_PRIME_BITS'd1199214675, `RNS_PRIME_BITS'd1878325668, `RNS_PRIME_BITS'd7727696, `RNS_PRIME_BITS'd909482893, `RNS_PRIME_BITS'd390894248, `RNS_PRIME_BITS'd791713145, `RNS_PRIME_BITS'd1215966900, `RNS_PRIME_BITS'd587075636, `RNS_PRIME_BITS'd1199234809, `RNS_PRIME_BITS'd39126152, `RNS_PRIME_BITS'd624524991, `RNS_PRIME_BITS'd1200643284, `RNS_PRIME_BITS'd2068724100, `RNS_PRIME_BITS'd1028019199, `RNS_PRIME_BITS'd764503116, `RNS_PRIME_BITS'd956844079, `RNS_PRIME_BITS'd976022455, `RNS_PRIME_BITS'd128768493, `RNS_PRIME_BITS'd601425161, `RNS_PRIME_BITS'd297804970, `RNS_PRIME_BITS'd86626384, `RNS_PRIME_BITS'd1057658604, `RNS_PRIME_BITS'd1158945815},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1180811958, `RNS_PRIME_BITS'd698897645, `RNS_PRIME_BITS'd396752410, `RNS_PRIME_BITS'd1590960824, `RNS_PRIME_BITS'd676858767, `RNS_PRIME_BITS'd1242864821, `RNS_PRIME_BITS'd1981568237, `RNS_PRIME_BITS'd2047801397, `RNS_PRIME_BITS'd1141109968, `RNS_PRIME_BITS'd640452388, `RNS_PRIME_BITS'd1735615176, `RNS_PRIME_BITS'd104371406, `RNS_PRIME_BITS'd793743842, `RNS_PRIME_BITS'd1404190271, `RNS_PRIME_BITS'd404036694, `RNS_PRIME_BITS'd2100155542, `RNS_PRIME_BITS'd1947317042, `RNS_PRIME_BITS'd1002584402, `RNS_PRIME_BITS'd1972104903, `RNS_PRIME_BITS'd1117302355, `RNS_PRIME_BITS'd1082672190, `RNS_PRIME_BITS'd665909595, `RNS_PRIME_BITS'd325883975, `RNS_PRIME_BITS'd1855667154, `RNS_PRIME_BITS'd536371151, `RNS_PRIME_BITS'd431097772, `RNS_PRIME_BITS'd1527060402, `RNS_PRIME_BITS'd1113343725, `RNS_PRIME_BITS'd1952670695, `RNS_PRIME_BITS'd1494908283, `RNS_PRIME_BITS'd1889283537, `RNS_PRIME_BITS'd524962442, `RNS_PRIME_BITS'd1401061297, `RNS_PRIME_BITS'd1349253646, `RNS_PRIME_BITS'd818503666, `RNS_PRIME_BITS'd723680490, `RNS_PRIME_BITS'd322476241, `RNS_PRIME_BITS'd1874038872, `RNS_PRIME_BITS'd834025286, `RNS_PRIME_BITS'd281055234, `RNS_PRIME_BITS'd1074140584, `RNS_PRIME_BITS'd49981851, `RNS_PRIME_BITS'd878592647, `RNS_PRIME_BITS'd1280361918, `RNS_PRIME_BITS'd1657938546, `RNS_PRIME_BITS'd658448763, `RNS_PRIME_BITS'd1234006662, `RNS_PRIME_BITS'd1800184525, `RNS_PRIME_BITS'd1599760116, `RNS_PRIME_BITS'd1944520926, `RNS_PRIME_BITS'd1201959893, `RNS_PRIME_BITS'd1601517741, `RNS_PRIME_BITS'd366288311, `RNS_PRIME_BITS'd1067917992, `RNS_PRIME_BITS'd1471009666, `RNS_PRIME_BITS'd1724844730, `RNS_PRIME_BITS'd1186389507, `RNS_PRIME_BITS'd1232517567, `RNS_PRIME_BITS'd2054892602, `RNS_PRIME_BITS'd1556827466, `RNS_PRIME_BITS'd971038417, `RNS_PRIME_BITS'd2023717671, `RNS_PRIME_BITS'd1674979427},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd863581131, `RNS_PRIME_BITS'd266488565, `RNS_PRIME_BITS'd197474481, `RNS_PRIME_BITS'd2131754249, `RNS_PRIME_BITS'd1844273609, `RNS_PRIME_BITS'd2052452190, `RNS_PRIME_BITS'd1532049341, `RNS_PRIME_BITS'd1811004807, `RNS_PRIME_BITS'd1970163605, `RNS_PRIME_BITS'd1802277828, `RNS_PRIME_BITS'd200129577, `RNS_PRIME_BITS'd1902288884, `RNS_PRIME_BITS'd600242329, `RNS_PRIME_BITS'd400413469, `RNS_PRIME_BITS'd735419640, `RNS_PRIME_BITS'd10234283, `RNS_PRIME_BITS'd1236975143, `RNS_PRIME_BITS'd354809650, `RNS_PRIME_BITS'd1260290827, `RNS_PRIME_BITS'd240751673, `RNS_PRIME_BITS'd2076469305, `RNS_PRIME_BITS'd231305546, `RNS_PRIME_BITS'd122535444, `RNS_PRIME_BITS'd1634152440, `RNS_PRIME_BITS'd449910378, `RNS_PRIME_BITS'd1239381293, `RNS_PRIME_BITS'd2113046598, `RNS_PRIME_BITS'd1065183214, `RNS_PRIME_BITS'd523000083, `RNS_PRIME_BITS'd831666628, `RNS_PRIME_BITS'd138524561, `RNS_PRIME_BITS'd1172437812, `RNS_PRIME_BITS'd590795774, `RNS_PRIME_BITS'd348980417, `RNS_PRIME_BITS'd1897963711, `RNS_PRIME_BITS'd1718005309, `RNS_PRIME_BITS'd1133296249, `RNS_PRIME_BITS'd796514801, `RNS_PRIME_BITS'd958676669, `RNS_PRIME_BITS'd64563004, `RNS_PRIME_BITS'd1975647812, `RNS_PRIME_BITS'd579138741, `RNS_PRIME_BITS'd36175035, `RNS_PRIME_BITS'd182951808, `RNS_PRIME_BITS'd1491813251, `RNS_PRIME_BITS'd1193767449, `RNS_PRIME_BITS'd1756567829, `RNS_PRIME_BITS'd1221476635, `RNS_PRIME_BITS'd1663696998, `RNS_PRIME_BITS'd1660937547, `RNS_PRIME_BITS'd19608843, `RNS_PRIME_BITS'd1804134098, `RNS_PRIME_BITS'd1143024219, `RNS_PRIME_BITS'd887687435, `RNS_PRIME_BITS'd1287398144, `RNS_PRIME_BITS'd120671020, `RNS_PRIME_BITS'd660093495, `RNS_PRIME_BITS'd1773444005, `RNS_PRIME_BITS'd960444154, `RNS_PRIME_BITS'd1827198507, `RNS_PRIME_BITS'd1783905120, `RNS_PRIME_BITS'd577134207, `RNS_PRIME_BITS'd708871736},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd2006888302, `RNS_PRIME_BITS'd1915797300, `RNS_PRIME_BITS'd49249814, `RNS_PRIME_BITS'd1610378484, `RNS_PRIME_BITS'd808269908, `RNS_PRIME_BITS'd1579153117, `RNS_PRIME_BITS'd785126063, `RNS_PRIME_BITS'd1519044505, `RNS_PRIME_BITS'd1343154438, `RNS_PRIME_BITS'd106304448, `RNS_PRIME_BITS'd1361590782, `RNS_PRIME_BITS'd408243051, `RNS_PRIME_BITS'd1624358720, `RNS_PRIME_BITS'd1076916254, `RNS_PRIME_BITS'd1411883997, `RNS_PRIME_BITS'd1499897549, `RNS_PRIME_BITS'd995275098, `RNS_PRIME_BITS'd573382855, `RNS_PRIME_BITS'd796043708, `RNS_PRIME_BITS'd1898906447, `RNS_PRIME_BITS'd2046261189, `RNS_PRIME_BITS'd1898694097, `RNS_PRIME_BITS'd1866665936, `RNS_PRIME_BITS'd321460536, `RNS_PRIME_BITS'd1935227906, `RNS_PRIME_BITS'd292174375, `RNS_PRIME_BITS'd1651256030, `RNS_PRIME_BITS'd1674111577, `RNS_PRIME_BITS'd362735615, `RNS_PRIME_BITS'd303641034, `RNS_PRIME_BITS'd136679130, `RNS_PRIME_BITS'd947974746, `RNS_PRIME_BITS'd1971088069, `RNS_PRIME_BITS'd331719264, `RNS_PRIME_BITS'd1067104690, `RNS_PRIME_BITS'd1014920853, `RNS_PRIME_BITS'd447649351, `RNS_PRIME_BITS'd305771017, `RNS_PRIME_BITS'd959695467, `RNS_PRIME_BITS'd731192465, `RNS_PRIME_BITS'd596300382, `RNS_PRIME_BITS'd1769119785, `RNS_PRIME_BITS'd1902426573, `RNS_PRIME_BITS'd654833583, `RNS_PRIME_BITS'd873629554, `RNS_PRIME_BITS'd711101770, `RNS_PRIME_BITS'd679149815, `RNS_PRIME_BITS'd558407411, `RNS_PRIME_BITS'd449470596, `RNS_PRIME_BITS'd276205002, `RNS_PRIME_BITS'd1788733215, `RNS_PRIME_BITS'd429865127, `RNS_PRIME_BITS'd1275811230, `RNS_PRIME_BITS'd1370277766, `RNS_PRIME_BITS'd1168169987, `RNS_PRIME_BITS'd538488167, `RNS_PRIME_BITS'd126138005, `RNS_PRIME_BITS'd1843645976, `RNS_PRIME_BITS'd342817420, `RNS_PRIME_BITS'd667896261, `RNS_PRIME_BITS'd1326718868, `RNS_PRIME_BITS'd1772889814, `RNS_PRIME_BITS'd1423092132},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd827630191, `RNS_PRIME_BITS'd634442553, `RNS_PRIME_BITS'd14124402, `RNS_PRIME_BITS'd1687474151, `RNS_PRIME_BITS'd14861374, `RNS_PRIME_BITS'd1248849378, `RNS_PRIME_BITS'd2105098028, `RNS_PRIME_BITS'd1655854283, `RNS_PRIME_BITS'd1376784415, `RNS_PRIME_BITS'd1875735111, `RNS_PRIME_BITS'd1629799445, `RNS_PRIME_BITS'd50859102, `RNS_PRIME_BITS'd353092123, `RNS_PRIME_BITS'd1463329648, `RNS_PRIME_BITS'd1971964208, `RNS_PRIME_BITS'd1351991644, `RNS_PRIME_BITS'd1423704554, `RNS_PRIME_BITS'd462906762, `RNS_PRIME_BITS'd1662891139, `RNS_PRIME_BITS'd1537383243, `RNS_PRIME_BITS'd190823532, `RNS_PRIME_BITS'd754518586, `RNS_PRIME_BITS'd1472669913, `RNS_PRIME_BITS'd1403908978, `RNS_PRIME_BITS'd838777520, `RNS_PRIME_BITS'd356624563, `RNS_PRIME_BITS'd1854365554, `RNS_PRIME_BITS'd1405622643, `RNS_PRIME_BITS'd182689866, `RNS_PRIME_BITS'd2088866633, `RNS_PRIME_BITS'd1993147357, `RNS_PRIME_BITS'd335862598, `RNS_PRIME_BITS'd520746293, `RNS_PRIME_BITS'd795266135, `RNS_PRIME_BITS'd276444971, `RNS_PRIME_BITS'd1008493454, `RNS_PRIME_BITS'd1962983607, `RNS_PRIME_BITS'd737870517, `RNS_PRIME_BITS'd140078324, `RNS_PRIME_BITS'd608663139, `RNS_PRIME_BITS'd481530671, `RNS_PRIME_BITS'd1794412482, `RNS_PRIME_BITS'd944136518, `RNS_PRIME_BITS'd1479984746, `RNS_PRIME_BITS'd1020523066, `RNS_PRIME_BITS'd1308174171, `RNS_PRIME_BITS'd129364822, `RNS_PRIME_BITS'd1843702908, `RNS_PRIME_BITS'd1806730708, `RNS_PRIME_BITS'd688071846, `RNS_PRIME_BITS'd2031608751, `RNS_PRIME_BITS'd1141675715, `RNS_PRIME_BITS'd2018762224, `RNS_PRIME_BITS'd999896244, `RNS_PRIME_BITS'd703901652, `RNS_PRIME_BITS'd1469183668, `RNS_PRIME_BITS'd1633319106, `RNS_PRIME_BITS'd541653944, `RNS_PRIME_BITS'd1165857483, `RNS_PRIME_BITS'd187415820, `RNS_PRIME_BITS'd1347391675, `RNS_PRIME_BITS'd1947813149, `RNS_PRIME_BITS'd1192713535},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1925970851, `RNS_PRIME_BITS'd207695132, `RNS_PRIME_BITS'd148848534, `RNS_PRIME_BITS'd1761745303, `RNS_PRIME_BITS'd1020094163, `RNS_PRIME_BITS'd1296504500, `RNS_PRIME_BITS'd1590156063, `RNS_PRIME_BITS'd1828920336, `RNS_PRIME_BITS'd1528595831, `RNS_PRIME_BITS'd1612223517, `RNS_PRIME_BITS'd1146443053, `RNS_PRIME_BITS'd822124619, `RNS_PRIME_BITS'd373441180, `RNS_PRIME_BITS'd1599886708, `RNS_PRIME_BITS'd1819024442, `RNS_PRIME_BITS'd1343916693, `RNS_PRIME_BITS'd1580226385, `RNS_PRIME_BITS'd1465397025, `RNS_PRIME_BITS'd576340174, `RNS_PRIME_BITS'd508007782, `RNS_PRIME_BITS'd1949278380, `RNS_PRIME_BITS'd1026065501, `RNS_PRIME_BITS'd1982388385, `RNS_PRIME_BITS'd601571399, `RNS_PRIME_BITS'd1814968618, `RNS_PRIME_BITS'd1139796275, `RNS_PRIME_BITS'd1376844757, `RNS_PRIME_BITS'd591326689, `RNS_PRIME_BITS'd284129690, `RNS_PRIME_BITS'd1468519535, `RNS_PRIME_BITS'd827950938, `RNS_PRIME_BITS'd1331495236, `RNS_PRIME_BITS'd1575358450, `RNS_PRIME_BITS'd368435717, `RNS_PRIME_BITS'd1380291710, `RNS_PRIME_BITS'd353025982, `RNS_PRIME_BITS'd228998489, `RNS_PRIME_BITS'd1188901935, `RNS_PRIME_BITS'd1389915387, `RNS_PRIME_BITS'd464898846, `RNS_PRIME_BITS'd1250107969, `RNS_PRIME_BITS'd622888137, `RNS_PRIME_BITS'd87729872, `RNS_PRIME_BITS'd1083576085, `RNS_PRIME_BITS'd1840014191, `RNS_PRIME_BITS'd1453536448, `RNS_PRIME_BITS'd1893528272, `RNS_PRIME_BITS'd824257829, `RNS_PRIME_BITS'd923463583, `RNS_PRIME_BITS'd1538410082, `RNS_PRIME_BITS'd1174453731, `RNS_PRIME_BITS'd911258653, `RNS_PRIME_BITS'd712118336, `RNS_PRIME_BITS'd1078820638, `RNS_PRIME_BITS'd1901471095, `RNS_PRIME_BITS'd768800080, `RNS_PRIME_BITS'd1427536931, `RNS_PRIME_BITS'd1721350193, `RNS_PRIME_BITS'd421031535, `RNS_PRIME_BITS'd1756461716, `RNS_PRIME_BITS'd1423546356, `RNS_PRIME_BITS'd181657083, `RNS_PRIME_BITS'd1451070185},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd679082962, `RNS_PRIME_BITS'd21725588, `RNS_PRIME_BITS'd1645223958, `RNS_PRIME_BITS'd1935386753, `RNS_PRIME_BITS'd147309818, `RNS_PRIME_BITS'd1358855180, `RNS_PRIME_BITS'd1309811091, `RNS_PRIME_BITS'd1178694670, `RNS_PRIME_BITS'd1626480704, `RNS_PRIME_BITS'd789699425, `RNS_PRIME_BITS'd1362151287, `RNS_PRIME_BITS'd1335637725, `RNS_PRIME_BITS'd799792040, `RNS_PRIME_BITS'd1787703015, `RNS_PRIME_BITS'd1889383441, `RNS_PRIME_BITS'd376392512, `RNS_PRIME_BITS'd1203126727, `RNS_PRIME_BITS'd649865995, `RNS_PRIME_BITS'd1898940369, `RNS_PRIME_BITS'd1306763942, `RNS_PRIME_BITS'd896631706, `RNS_PRIME_BITS'd1233985319, `RNS_PRIME_BITS'd1297846148, `RNS_PRIME_BITS'd1971934677, `RNS_PRIME_BITS'd1424335466, `RNS_PRIME_BITS'd216329546, `RNS_PRIME_BITS'd1938315192, `RNS_PRIME_BITS'd1163148101, `RNS_PRIME_BITS'd1843731486, `RNS_PRIME_BITS'd2000376334, `RNS_PRIME_BITS'd153601635, `RNS_PRIME_BITS'd1410137926, `RNS_PRIME_BITS'd476307234, `RNS_PRIME_BITS'd489843704, `RNS_PRIME_BITS'd1154289721, `RNS_PRIME_BITS'd741963136, `RNS_PRIME_BITS'd205108911, `RNS_PRIME_BITS'd1051329728, `RNS_PRIME_BITS'd881212437, `RNS_PRIME_BITS'd1454002446, `RNS_PRIME_BITS'd59717368, `RNS_PRIME_BITS'd1546369699, `RNS_PRIME_BITS'd1009475440, `RNS_PRIME_BITS'd539509008, `RNS_PRIME_BITS'd341138130, `RNS_PRIME_BITS'd1720619438, `RNS_PRIME_BITS'd535596838, `RNS_PRIME_BITS'd1631833303, `RNS_PRIME_BITS'd933766656, `RNS_PRIME_BITS'd926729148, `RNS_PRIME_BITS'd1837590264, `RNS_PRIME_BITS'd621781956, `RNS_PRIME_BITS'd2122931229, `RNS_PRIME_BITS'd2098610929, `RNS_PRIME_BITS'd863275331, `RNS_PRIME_BITS'd1075515373, `RNS_PRIME_BITS'd375638505, `RNS_PRIME_BITS'd665726026, `RNS_PRIME_BITS'd467316107, `RNS_PRIME_BITS'd547754318, `RNS_PRIME_BITS'd1580566206, `RNS_PRIME_BITS'd802589102, `RNS_PRIME_BITS'd148205767},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd985627742, `RNS_PRIME_BITS'd209219715, `RNS_PRIME_BITS'd1797297359, `RNS_PRIME_BITS'd607947504, `RNS_PRIME_BITS'd582137866, `RNS_PRIME_BITS'd1553772574, `RNS_PRIME_BITS'd1001224375, `RNS_PRIME_BITS'd408115440, `RNS_PRIME_BITS'd1688164042, `RNS_PRIME_BITS'd1138957206, `RNS_PRIME_BITS'd29488642, `RNS_PRIME_BITS'd695959640, `RNS_PRIME_BITS'd1479303328, `RNS_PRIME_BITS'd519154132, `RNS_PRIME_BITS'd963399678, `RNS_PRIME_BITS'd405602459, `RNS_PRIME_BITS'd1892086515, `RNS_PRIME_BITS'd80644722, `RNS_PRIME_BITS'd1766908121, `RNS_PRIME_BITS'd589212064, `RNS_PRIME_BITS'd1938421324, `RNS_PRIME_BITS'd223488580, `RNS_PRIME_BITS'd1007863781, `RNS_PRIME_BITS'd572067441, `RNS_PRIME_BITS'd1628177047, `RNS_PRIME_BITS'd70232036, `RNS_PRIME_BITS'd888471290, `RNS_PRIME_BITS'd41854895, `RNS_PRIME_BITS'd369428266, `RNS_PRIME_BITS'd980564471, `RNS_PRIME_BITS'd1490691155, `RNS_PRIME_BITS'd37028611, `RNS_PRIME_BITS'd2016849603, `RNS_PRIME_BITS'd269448364, `RNS_PRIME_BITS'd1080531861, `RNS_PRIME_BITS'd117506787, `RNS_PRIME_BITS'd1446317206, `RNS_PRIME_BITS'd1362925816, `RNS_PRIME_BITS'd702116429, `RNS_PRIME_BITS'd1232945780, `RNS_PRIME_BITS'd410918689, `RNS_PRIME_BITS'd156420353, `RNS_PRIME_BITS'd901760470, `RNS_PRIME_BITS'd1589572379, `RNS_PRIME_BITS'd472182866, `RNS_PRIME_BITS'd1578477615, `RNS_PRIME_BITS'd1370829515, `RNS_PRIME_BITS'd2028194232, `RNS_PRIME_BITS'd971006858, `RNS_PRIME_BITS'd908554640, `RNS_PRIME_BITS'd768568972, `RNS_PRIME_BITS'd202469597, `RNS_PRIME_BITS'd1343706043, `RNS_PRIME_BITS'd387366877, `RNS_PRIME_BITS'd1612097702, `RNS_PRIME_BITS'd316054804, `RNS_PRIME_BITS'd400914411, `RNS_PRIME_BITS'd828730173, `RNS_PRIME_BITS'd786533504, `RNS_PRIME_BITS'd574179569, `RNS_PRIME_BITS'd935110882, `RNS_PRIME_BITS'd796989334, `RNS_PRIME_BITS'd732343142}
};
parameter q_BASIS_poly untwist_factor_q = '{
    '{`RNS_PRIME_BITS'd253, `RNS_PRIME_BITS'd228, `RNS_PRIME_BITS'd111, `RNS_PRIME_BITS'd98, `RNS_PRIME_BITS'd68, `RNS_PRIME_BITS'd236, `RNS_PRIME_BITS'd169, `RNS_PRIME_BITS'd133, `RNS_PRIME_BITS'd129, `RNS_PRIME_BITS'd100, `RNS_PRIME_BITS'd211, `RNS_PRIME_BITS'd52, `RNS_PRIME_BITS'd120, `RNS_PRIME_BITS'd99, `RNS_PRIME_BITS'd11, `RNS_PRIME_BITS'd144, `RNS_PRIME_BITS'd16, `RNS_PRIME_BITS'd116, `RNS_PRIME_BITS'd70, `RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd242, `RNS_PRIME_BITS'd84, `RNS_PRIME_BITS'd95, `RNS_PRIME_BITS'd239, `RNS_PRIME_BITS'd255, `RNS_PRIME_BITS'd114, `RNS_PRIME_BITS'd184, `RNS_PRIME_BITS'd49, `RNS_PRIME_BITS'd34, `RNS_PRIME_BITS'd118, `RNS_PRIME_BITS'd213, `RNS_PRIME_BITS'd195, `RNS_PRIME_BITS'd193, `RNS_PRIME_BITS'd50, `RNS_PRIME_BITS'd234, `RNS_PRIME_BITS'd26, `RNS_PRIME_BITS'd60, `RNS_PRIME_BITS'd178, `RNS_PRIME_BITS'd134, `RNS_PRIME_BITS'd72, `RNS_PRIME_BITS'd8, `RNS_PRIME_BITS'd58, `RNS_PRIME_BITS'd35, `RNS_PRIME_BITS'd61, `RNS_PRIME_BITS'd121, `RNS_PRIME_BITS'd42, `RNS_PRIME_BITS'd176, `RNS_PRIME_BITS'd248, `RNS_PRIME_BITS'd256, `RNS_PRIME_BITS'd57, `RNS_PRIME_BITS'd92, `RNS_PRIME_BITS'd153, `RNS_PRIME_BITS'd17, `RNS_PRIME_BITS'd59, `RNS_PRIME_BITS'd235, `RNS_PRIME_BITS'd226, `RNS_PRIME_BITS'd225, `RNS_PRIME_BITS'd25, `RNS_PRIME_BITS'd117, `RNS_PRIME_BITS'd13, `RNS_PRIME_BITS'd30, `RNS_PRIME_BITS'd89, `RNS_PRIME_BITS'd67, `RNS_PRIME_BITS'd36},
    '{`RNS_PRIME_BITS'd2113929343, `RNS_PRIME_BITS'd719749060, `RNS_PRIME_BITS'd1215239054, `RNS_PRIME_BITS'd1721455720, `RNS_PRIME_BITS'd1048303337, `RNS_PRIME_BITS'd265552380, `RNS_PRIME_BITS'd1471263777, `RNS_PRIME_BITS'd600370338, `RNS_PRIME_BITS'd1711251046, `RNS_PRIME_BITS'd1039522340, `RNS_PRIME_BITS'd969189398, `RNS_PRIME_BITS'd83871020, `RNS_PRIME_BITS'd34507746, `RNS_PRIME_BITS'd699166695, `RNS_PRIME_BITS'd1390803476, `RNS_PRIME_BITS'd1022064446, `RNS_PRIME_BITS'd254214852, `RNS_PRIME_BITS'd1301117692, `RNS_PRIME_BITS'd1833562202, `RNS_PRIME_BITS'd584132787, `RNS_PRIME_BITS'd875293636, `RNS_PRIME_BITS'd17774605, `RNS_PRIME_BITS'd356785962, `RNS_PRIME_BITS'd2038988113, `RNS_PRIME_BITS'd955160690, `RNS_PRIME_BITS'd1328378368, `RNS_PRIME_BITS'd1144173285, `RNS_PRIME_BITS'd781130222, `RNS_PRIME_BITS'd268845809, `RNS_PRIME_BITS'd1825799892, `RNS_PRIME_BITS'd1240852021, `RNS_PRIME_BITS'd1464300718, `RNS_PRIME_BITS'd386689036, `RNS_PRIME_BITS'd1486183251, `RNS_PRIME_BITS'd1368379953, `RNS_PRIME_BITS'd1119124109, `RNS_PRIME_BITS'd1748752439, `RNS_PRIME_BITS'd957539307, `RNS_PRIME_BITS'd1125311264, `RNS_PRIME_BITS'd2055724711, `RNS_PRIME_BITS'd1973052422, `RNS_PRIME_BITS'd626565169, `RNS_PRIME_BITS'd713461989, `RNS_PRIME_BITS'd33303951, `RNS_PRIME_BITS'd350105513, `RNS_PRIME_BITS'd1455447908, `RNS_PRIME_BITS'd1831138265, `RNS_PRIME_BITS'd1405399662, `RNS_PRIME_BITS'd184742794, `RNS_PRIME_BITS'd1044496195, `RNS_PRIME_BITS'd761311156, `RNS_PRIME_BITS'd1053061321, `RNS_PRIME_BITS'd1242777573, `RNS_PRIME_BITS'd519640201, `RNS_PRIME_BITS'd1978003332, `RNS_PRIME_BITS'd1147003102, `RNS_PRIME_BITS'd12870039, `RNS_PRIME_BITS'd1358866390, `RNS_PRIME_BITS'd694384824, `RNS_PRIME_BITS'd967763240, `RNS_PRIME_BITS'd1675838128, `RNS_PRIME_BITS'd1614885743, `RNS_PRIME_BITS'd577663718, `RNS_PRIME_BITS'd1655002074},
    '{`RNS_PRIME_BITS'd2113929721, `RNS_PRIME_BITS'd1129628573, `RNS_PRIME_BITS'd1261982508, `RNS_PRIME_BITS'd1269054906, `RNS_PRIME_BITS'd2006306856, `RNS_PRIME_BITS'd1549546859, `RNS_PRIME_BITS'd2055709882, `RNS_PRIME_BITS'd2108038524, `RNS_PRIME_BITS'd1738613598, `RNS_PRIME_BITS'd171013086, `RNS_PRIME_BITS'd1930778971, `RNS_PRIME_BITS'd768892011, `RNS_PRIME_BITS'd670592079, `RNS_PRIME_BITS'd801729623, `RNS_PRIME_BITS'd333776617, `RNS_PRIME_BITS'd643203401, `RNS_PRIME_BITS'd1056112510, `RNS_PRIME_BITS'd121712876, `RNS_PRIME_BITS'd1086361181, `RNS_PRIME_BITS'd695697577, `RNS_PRIME_BITS'd2051130920, `RNS_PRIME_BITS'd344670759, `RNS_PRIME_BITS'd848493897, `RNS_PRIME_BITS'd611046607, `RNS_PRIME_BITS'd2011563958, `RNS_PRIME_BITS'd1065701949, `RNS_PRIME_BITS'd335008896, `RNS_PRIME_BITS'd1566302183, `RNS_PRIME_BITS'd816075104, `RNS_PRIME_BITS'd247813306, `RNS_PRIME_BITS'd1799236445, `RNS_PRIME_BITS'd158825453, `RNS_PRIME_BITS'd1972921725, `RNS_PRIME_BITS'd692318239, `RNS_PRIME_BITS'd281004805, `RNS_PRIME_BITS'd141147247, `RNS_PRIME_BITS'd581229285, `RNS_PRIME_BITS'd1386640185, `RNS_PRIME_BITS'd389570102, `RNS_PRIME_BITS'd1152721697, `RNS_PRIME_BITS'd2050935508, `RNS_PRIME_BITS'd678148867, `RNS_PRIME_BITS'd2071007759, `RNS_PRIME_BITS'd251669112, `RNS_PRIME_BITS'd961135379, `RNS_PRIME_BITS'd1972902860, `RNS_PRIME_BITS'd1676556220, `RNS_PRIME_BITS'd1009669518, `RNS_PRIME_BITS'd336386816, `RNS_PRIME_BITS'd151883032, `RNS_PRIME_BITS'd774727052, `RNS_PRIME_BITS'd1242808425, `RNS_PRIME_BITS'd1480771520, `RNS_PRIME_BITS'd944885152, `RNS_PRIME_BITS'd478263574, `RNS_PRIME_BITS'd221482402, `RNS_PRIME_BITS'd278774359, `RNS_PRIME_BITS'd1534498320, `RNS_PRIME_BITS'd2033364169, `RNS_PRIME_BITS'd1427971716, `RNS_PRIME_BITS'd468707300, `RNS_PRIME_BITS'd1859106025, `RNS_PRIME_BITS'd1235052902, `RNS_PRIME_BITS'd1377669667},
    '{`RNS_PRIME_BITS'd2113930477, `RNS_PRIME_BITS'd753643868, `RNS_PRIME_BITS'd1459869973, `RNS_PRIME_BITS'd535517695, `RNS_PRIME_BITS'd1404633782, `RNS_PRIME_BITS'd292592800, `RNS_PRIME_BITS'd1507938333, `RNS_PRIME_BITS'd1830244510, `RNS_PRIME_BITS'd1562108556, `RNS_PRIME_BITS'd390708063, `RNS_PRIME_BITS'd2097867677, `RNS_PRIME_BITS'd101893994, `RNS_PRIME_BITS'd652328989, `RNS_PRIME_BITS'd2104172274, `RNS_PRIME_BITS'd267824270, `RNS_PRIME_BITS'd1893865721, `RNS_PRIME_BITS'd1735658448, `RNS_PRIME_BITS'd1725832022, `RNS_PRIME_BITS'd1900233247, `RNS_PRIME_BITS'd1336070358, `RNS_PRIME_BITS'd421997206, `RNS_PRIME_BITS'd536750487, `RNS_PRIME_BITS'd1178611434, `RNS_PRIME_BITS'd618796859, `RNS_PRIME_BITS'd1472788446, `RNS_PRIME_BITS'd2121645181, `RNS_PRIME_BITS'd1491675868, `RNS_PRIME_BITS'd2003607145, `RNS_PRIME_BITS'd934272159, `RNS_PRIME_BITS'd225220907, `RNS_PRIME_BITS'd480194134, `RNS_PRIME_BITS'd48193229, `RNS_PRIME_BITS'd1751633961, `RNS_PRIME_BITS'd1708385398, `RNS_PRIME_BITS'd29758940, `RNS_PRIME_BITS'd1977645907, `RNS_PRIME_BITS'd756157563, `RNS_PRIME_BITS'd264416368, `RNS_PRIME_BITS'd830221424, `RNS_PRIME_BITS'd1920620573, `RNS_PRIME_BITS'd1199928760, `RNS_PRIME_BITS'd1413085432, `RNS_PRIME_BITS'd1074126258, `RNS_PRIME_BITS'd871527458, `RNS_PRIME_BITS'd1546300093, `RNS_PRIME_BITS'd718563074, `RNS_PRIME_BITS'd2126107401, `RNS_PRIME_BITS'd423807776, `RNS_PRIME_BITS'd633795346, `RNS_PRIME_BITS'd90794750, `RNS_PRIME_BITS'd1195992423, `RNS_PRIME_BITS'd1686683653, `RNS_PRIME_BITS'd655871583, `RNS_PRIME_BITS'd970106672, `RNS_PRIME_BITS'd1785392179, `RNS_PRIME_BITS'd1824474512, `RNS_PRIME_BITS'd999290885, `RNS_PRIME_BITS'd108997519, `RNS_PRIME_BITS'd453130443, `RNS_PRIME_BITS'd494910485, `RNS_PRIME_BITS'd799885904, `RNS_PRIME_BITS'd625570152, `RNS_PRIME_BITS'd1798892458, `RNS_PRIME_BITS'd1984677102},
    '{`RNS_PRIME_BITS'd2113930603, `RNS_PRIME_BITS'd1148234337, `RNS_PRIME_BITS'd1277003118, `RNS_PRIME_BITS'd555253243, `RNS_PRIME_BITS'd311219111, `RNS_PRIME_BITS'd1914050636, `RNS_PRIME_BITS'd2094672516, `RNS_PRIME_BITS'd82126026, `RNS_PRIME_BITS'd1919207634, `RNS_PRIME_BITS'd44124382, `RNS_PRIME_BITS'd1325491942, `RNS_PRIME_BITS'd1839771716, `RNS_PRIME_BITS'd1484926716, `RNS_PRIME_BITS'd685862911, `RNS_PRIME_BITS'd976250481, `RNS_PRIME_BITS'd1719835357, `RNS_PRIME_BITS'd408080019, `RNS_PRIME_BITS'd182045370, `RNS_PRIME_BITS'd1969424525, `RNS_PRIME_BITS'd1651817411, `RNS_PRIME_BITS'd2060370494, `RNS_PRIME_BITS'd221153168, `RNS_PRIME_BITS'd905189292, `RNS_PRIME_BITS'd1325394714, `RNS_PRIME_BITS'd62717420, `RNS_PRIME_BITS'd188295079, `RNS_PRIME_BITS'd776025039, `RNS_PRIME_BITS'd565387027, `RNS_PRIME_BITS'd1397979561, `RNS_PRIME_BITS'd1664933581, `RNS_PRIME_BITS'd448680268, `RNS_PRIME_BITS'd1622276664, `RNS_PRIME_BITS'd327342002, `RNS_PRIME_BITS'd540905663, `RNS_PRIME_BITS'd1956354845, `RNS_PRIME_BITS'd1278113227, `RNS_PRIME_BITS'd1492554435, `RNS_PRIME_BITS'd1653862382, `RNS_PRIME_BITS'd1469660074, `RNS_PRIME_BITS'd494936011, `RNS_PRIME_BITS'd574985373, `RNS_PRIME_BITS'd229789241, `RNS_PRIME_BITS'd895565421, `RNS_PRIME_BITS'd2063459396, `RNS_PRIME_BITS'd620076777, `RNS_PRIME_BITS'd204067039, `RNS_PRIME_BITS'd588314791, `RNS_PRIME_BITS'd1647295872, `RNS_PRIME_BITS'd705383058, `RNS_PRIME_BITS'd731884915, `RNS_PRIME_BITS'd2091990130, `RNS_PRIME_BITS'd1128449189, `RNS_PRIME_BITS'd468131553, `RNS_PRIME_BITS'd241316645, `RNS_PRIME_BITS'd1197953276, `RNS_PRIME_BITS'd519041421, `RNS_PRIME_BITS'd1746389166, `RNS_PRIME_BITS'd1478988427, `RNS_PRIME_BITS'd1758966300, `RNS_PRIME_BITS'd492740892, `RNS_PRIME_BITS'd1854190662, `RNS_PRIME_BITS'd866216548, `RNS_PRIME_BITS'd1499030155, `RNS_PRIME_BITS'd1793490330},
    '{`RNS_PRIME_BITS'd2113932367, `RNS_PRIME_BITS'd1867974872, `RNS_PRIME_BITS'd2104914645, `RNS_PRIME_BITS'd1045869907, `RNS_PRIME_BITS'd1414292750, `RNS_PRIME_BITS'd1931153017, `RNS_PRIME_BITS'd1213805772, `RNS_PRIME_BITS'd1835182550, `RNS_PRIME_BITS'd1474511724, `RNS_PRIME_BITS'd2127371253, `RNS_PRIME_BITS'd355229186, `RNS_PRIME_BITS'd888111261, `RNS_PRIME_BITS'd575791081, `RNS_PRIME_BITS'd368792914, `RNS_PRIME_BITS'd343147153, `RNS_PRIME_BITS'd1249075051, `RNS_PRIME_BITS'd886885442, `RNS_PRIME_BITS'd677197750, `RNS_PRIME_BITS'd820209434, `RNS_PRIME_BITS'd77353864, `RNS_PRIME_BITS'd2144628227, `RNS_PRIME_BITS'd1979149204, `RNS_PRIME_BITS'd1769338504, `RNS_PRIME_BITS'd103348431, `RNS_PRIME_BITS'd2012260124, `RNS_PRIME_BITS'd2031844080, `RNS_PRIME_BITS'd1631724075, `RNS_PRIME_BITS'd1894897721, `RNS_PRIME_BITS'd2019979570, `RNS_PRIME_BITS'd2084276684, `RNS_PRIME_BITS'd28101663, `RNS_PRIME_BITS'd2071146701, `RNS_PRIME_BITS'd1726513724, `RNS_PRIME_BITS'd568261748, `RNS_PRIME_BITS'd121223137, `RNS_PRIME_BITS'd629363282, `RNS_PRIME_BITS'd1526862685, `RNS_PRIME_BITS'd168310539, `RNS_PRIME_BITS'd1490586358, `RNS_PRIME_BITS'd1402258395, `RNS_PRIME_BITS'd1853517361, `RNS_PRIME_BITS'd669175024, `RNS_PRIME_BITS'd331930671, `RNS_PRIME_BITS'd1880160642, `RNS_PRIME_BITS'd1908843730, `RNS_PRIME_BITS'd349407258, `RNS_PRIME_BITS'd1672180200, `RNS_PRIME_BITS'd1289297062, `RNS_PRIME_BITS'd1442682816, `RNS_PRIME_BITS'd1867560061, `RNS_PRIME_BITS'd966823518, `RNS_PRIME_BITS'd829483264, `RNS_PRIME_BITS'd1715109801, `RNS_PRIME_BITS'd1372606738, `RNS_PRIME_BITS'd106057337, `RNS_PRIME_BITS'd673860316, `RNS_PRIME_BITS'd206584424, `RNS_PRIME_BITS'd2022885132, `RNS_PRIME_BITS'd974564895, `RNS_PRIME_BITS'd273173563, `RNS_PRIME_BITS'd268681678, `RNS_PRIME_BITS'd1641084080, `RNS_PRIME_BITS'd1774223663, `RNS_PRIME_BITS'd355605847},
    '{`RNS_PRIME_BITS'd2113933501, `RNS_PRIME_BITS'd1185726186, `RNS_PRIME_BITS'd710497597, `RNS_PRIME_BITS'd650360018, `RNS_PRIME_BITS'd157336621, `RNS_PRIME_BITS'd397297478, `RNS_PRIME_BITS'd776501032, `RNS_PRIME_BITS'd702673594, `RNS_PRIME_BITS'd1300211623, `RNS_PRIME_BITS'd82410844, `RNS_PRIME_BITS'd179916410, `RNS_PRIME_BITS'd986700450, `RNS_PRIME_BITS'd1301908858, `RNS_PRIME_BITS'd1012240544, `RNS_PRIME_BITS'd331229297, `RNS_PRIME_BITS'd127195022, `RNS_PRIME_BITS'd1702554385, `RNS_PRIME_BITS'd1834885785, `RNS_PRIME_BITS'd324434035, `RNS_PRIME_BITS'd1664074539, `RNS_PRIME_BITS'd1566829726, `RNS_PRIME_BITS'd406483085, `RNS_PRIME_BITS'd1348092004, `RNS_PRIME_BITS'd997317807, `RNS_PRIME_BITS'd559001618, `RNS_PRIME_BITS'd1427848259, `RNS_PRIME_BITS'd297212828, `RNS_PRIME_BITS'd227886979, `RNS_PRIME_BITS'd688786362, `RNS_PRIME_BITS'd1661051490, `RNS_PRIME_BITS'd1068560887, `RNS_PRIME_BITS'd136974249, `RNS_PRIME_BITS'd857604895, `RNS_PRIME_BITS'd870281389, `RNS_PRIME_BITS'd330800609, `RNS_PRIME_BITS'd2108265757, `RNS_PRIME_BITS'd812704507, `RNS_PRIME_BITS'd980834125, `RNS_PRIME_BITS'd1304060276, `RNS_PRIME_BITS'd36871064, `RNS_PRIME_BITS'd1874029180, `RNS_PRIME_BITS'd507705345, `RNS_PRIME_BITS'd540759405, `RNS_PRIME_BITS'd135799669, `RNS_PRIME_BITS'd473647087, `RNS_PRIME_BITS'd2000831818, `RNS_PRIME_BITS'd225922393, `RNS_PRIME_BITS'd856865827, `RNS_PRIME_BITS'd412772601, `RNS_PRIME_BITS'd951019813, `RNS_PRIME_BITS'd989808184, `RNS_PRIME_BITS'd2122107396, `RNS_PRIME_BITS'd1436464703, `RNS_PRIME_BITS'd2059104145, `RNS_PRIME_BITS'd2145826994, `RNS_PRIME_BITS'd180340212, `RNS_PRIME_BITS'd815127430, `RNS_PRIME_BITS'd1564793906, `RNS_PRIME_BITS'd948406233, `RNS_PRIME_BITS'd658460783, `RNS_PRIME_BITS'd1719671837, `RNS_PRIME_BITS'd737429472, `RNS_PRIME_BITS'd1714899668, `RNS_PRIME_BITS'd1512149371},
    '{`RNS_PRIME_BITS'd2113935013, `RNS_PRIME_BITS'd2095298864, `RNS_PRIME_BITS'd942646616, `RNS_PRIME_BITS'd1958663922, `RNS_PRIME_BITS'd399725916, `RNS_PRIME_BITS'd350883241, `RNS_PRIME_BITS'd1870590002, `RNS_PRIME_BITS'd41588437, `RNS_PRIME_BITS'd1721879254, `RNS_PRIME_BITS'd660092017, `RNS_PRIME_BITS'd1729211870, `RNS_PRIME_BITS'd1579073993, `RNS_PRIME_BITS'd82824889, `RNS_PRIME_BITS'd1545318742, `RNS_PRIME_BITS'd1264320790, `RNS_PRIME_BITS'd642860313, `RNS_PRIME_BITS'd1984463583, `RNS_PRIME_BITS'd736178203, `RNS_PRIME_BITS'd885531927, `RNS_PRIME_BITS'd1930216720, `RNS_PRIME_BITS'd1386165247, `RNS_PRIME_BITS'd186575011, `RNS_PRIME_BITS'd39071353, `RNS_PRIME_BITS'd1569538712, `RNS_PRIME_BITS'd1164897979, `RNS_PRIME_BITS'd1742646525, `RNS_PRIME_BITS'd1766860546, `RNS_PRIME_BITS'd1814827202, `RNS_PRIME_BITS'd454005626, `RNS_PRIME_BITS'd1438525080, `RNS_PRIME_BITS'd759328019, `RNS_PRIME_BITS'd1770253112, `RNS_PRIME_BITS'd196079291, `RNS_PRIME_BITS'd941938269, `RNS_PRIME_BITS'd269352175, `RNS_PRIME_BITS'd332690711, `RNS_PRIME_BITS'd1689317871, `RNS_PRIME_BITS'd1648751739, `RNS_PRIME_BITS'd1705708466, `RNS_PRIME_BITS'd1597511254, `RNS_PRIME_BITS'd1655790123, `RNS_PRIME_BITS'd815852633, `RNS_PRIME_BITS'd1934373040, `RNS_PRIME_BITS'd1473417439, `RNS_PRIME_BITS'd345078151, `RNS_PRIME_BITS'd74680898, `RNS_PRIME_BITS'd328312322, `RNS_PRIME_BITS'd1387044625, `RNS_PRIME_BITS'd918401803, `RNS_PRIME_BITS'd1579805212, `RNS_PRIME_BITS'd1587752627, `RNS_PRIME_BITS'd900455084, `RNS_PRIME_BITS'd1005841047, `RNS_PRIME_BITS'd679179388, `RNS_PRIME_BITS'd205573307, `RNS_PRIME_BITS'd1018677988, `RNS_PRIME_BITS'd343227041, `RNS_PRIME_BITS'd1443506900, `RNS_PRIME_BITS'd1121340545, `RNS_PRIME_BITS'd2080148280, `RNS_PRIME_BITS'd1282259653, `RNS_PRIME_BITS'd1677505507, `RNS_PRIME_BITS'd1902694704, `RNS_PRIME_BITS'd1564130907},
    '{`RNS_PRIME_BITS'd2113936147, `RNS_PRIME_BITS'd1353063251, `RNS_PRIME_BITS'd1976879587, `RNS_PRIME_BITS'd1722593273, `RNS_PRIME_BITS'd643646126, `RNS_PRIME_BITS'd1570484857, `RNS_PRIME_BITS'd1617276462, `RNS_PRIME_BITS'd1152103706, `RNS_PRIME_BITS'd524860171, `RNS_PRIME_BITS'd1815789325, `RNS_PRIME_BITS'd989779688, `RNS_PRIME_BITS'd2136363840, `RNS_PRIME_BITS'd958843302, `RNS_PRIME_BITS'd1156058131, `RNS_PRIME_BITS'd1116816771, `RNS_PRIME_BITS'd1025761684, `RNS_PRIME_BITS'd1228639026, `RNS_PRIME_BITS'd507286293, `RNS_PRIME_BITS'd2124779182, `RNS_PRIME_BITS'd1548313253, `RNS_PRIME_BITS'd687714506, `RNS_PRIME_BITS'd535501893, `RNS_PRIME_BITS'd292258251, `RNS_PRIME_BITS'd14021605, `RNS_PRIME_BITS'd999372216, `RNS_PRIME_BITS'd1958000551, `RNS_PRIME_BITS'd1558486882, `RNS_PRIME_BITS'd835285449, `RNS_PRIME_BITS'd2074865574, `RNS_PRIME_BITS'd2058814547, `RNS_PRIME_BITS'd162015902, `RNS_PRIME_BITS'd1653112125, `RNS_PRIME_BITS'd113413555, `RNS_PRIME_BITS'd859481359, `RNS_PRIME_BITS'd1554117857, `RNS_PRIME_BITS'd867978566, `RNS_PRIME_BITS'd1098060407, `RNS_PRIME_BITS'd683132183, `RNS_PRIME_BITS'd1693472326, `RNS_PRIME_BITS'd1380931880, `RNS_PRIME_BITS'd225482241, `RNS_PRIME_BITS'd1076325068, `RNS_PRIME_BITS'd957049445, `RNS_PRIME_BITS'd1445942374, `RNS_PRIME_BITS'd1267134975, `RNS_PRIME_BITS'd460758273, `RNS_PRIME_BITS'd1084403058, `RNS_PRIME_BITS'd545736177, `RNS_PRIME_BITS'd683646684, `RNS_PRIME_BITS'd1917741180, `RNS_PRIME_BITS'd1719837955, `RNS_PRIME_BITS'd933692158, `RNS_PRIME_BITS'd356254265, `RNS_PRIME_BITS'd1492041218, `RNS_PRIME_BITS'd947890726, `RNS_PRIME_BITS'd1821615501, `RNS_PRIME_BITS'd508295792, `RNS_PRIME_BITS'd1015344614, `RNS_PRIME_BITS'd1724578302, `RNS_PRIME_BITS'd621597327, `RNS_PRIME_BITS'd744227196, `RNS_PRIME_BITS'd735874166, `RNS_PRIME_BITS'd936281940, `RNS_PRIME_BITS'd1144315676},
    '{`RNS_PRIME_BITS'd2113936651, `RNS_PRIME_BITS'd232566135, `RNS_PRIME_BITS'd1530968846, `RNS_PRIME_BITS'd2055685754, `RNS_PRIME_BITS'd461205039, `RNS_PRIME_BITS'd361798236, `RNS_PRIME_BITS'd325143531, `RNS_PRIME_BITS'd1369867199, `RNS_PRIME_BITS'd1493149823, `RNS_PRIME_BITS'd87174973, `RNS_PRIME_BITS'd1611382155, `RNS_PRIME_BITS'd939911150, `RNS_PRIME_BITS'd124502857, `RNS_PRIME_BITS'd1850342453, `RNS_PRIME_BITS'd1998792858, `RNS_PRIME_BITS'd2132901097, `RNS_PRIME_BITS'd746257255, `RNS_PRIME_BITS'd1266704200, `RNS_PRIME_BITS'd1516624622, `RNS_PRIME_BITS'd598651617, `RNS_PRIME_BITS'd528442972, `RNS_PRIME_BITS'd1594845347, `RNS_PRIME_BITS'd1150247224, `RNS_PRIME_BITS'd1878121717, `RNS_PRIME_BITS'd447044912, `RNS_PRIME_BITS'd690876606, `RNS_PRIME_BITS'd2131064174, `RNS_PRIME_BITS'd1573859024, `RNS_PRIME_BITS'd2135898027, `RNS_PRIME_BITS'd1894573574, `RNS_PRIME_BITS'd1871400993, `RNS_PRIME_BITS'd1133412400, `RNS_PRIME_BITS'd179293895, `RNS_PRIME_BITS'd1172009225, `RNS_PRIME_BITS'd438507820, `RNS_PRIME_BITS'd977828196, `RNS_PRIME_BITS'd149598561, `RNS_PRIME_BITS'd1848768626, `RNS_PRIME_BITS'd332165351, `RNS_PRIME_BITS'd1387035859, `RNS_PRIME_BITS'd673834071, `RNS_PRIME_BITS'd113939354, `RNS_PRIME_BITS'd1289346430, `RNS_PRIME_BITS'd858408430, `RNS_PRIME_BITS'd1254654714, `RNS_PRIME_BITS'd540756407, `RNS_PRIME_BITS'd358945894, `RNS_PRIME_BITS'd216082995, `RNS_PRIME_BITS'd2141610068, `RNS_PRIME_BITS'd540905734, `RNS_PRIME_BITS'd1280694591, `RNS_PRIME_BITS'd1329685250, `RNS_PRIME_BITS'd952212611, `RNS_PRIME_BITS'd1824216637, `RNS_PRIME_BITS'd1094961097, `RNS_PRIME_BITS'd2122077440, `RNS_PRIME_BITS'd451346596, `RNS_PRIME_BITS'd617070652, `RNS_PRIME_BITS'd381422488, `RNS_PRIME_BITS'd1943862185, `RNS_PRIME_BITS'd3314132, `RNS_PRIME_BITS'd712493476, `RNS_PRIME_BITS'd670751538, `RNS_PRIME_BITS'd593371229},
    '{`RNS_PRIME_BITS'd2113937785, `RNS_PRIME_BITS'd1263630723, `RNS_PRIME_BITS'd725747538, `RNS_PRIME_BITS'd1126244205, `RNS_PRIME_BITS'd1635202277, `RNS_PRIME_BITS'd2135202767, `RNS_PRIME_BITS'd2033879740, `RNS_PRIME_BITS'd1436582137, `RNS_PRIME_BITS'd666153004, `RNS_PRIME_BITS'd1249884558, `RNS_PRIME_BITS'd967029865, `RNS_PRIME_BITS'd1958724106, `RNS_PRIME_BITS'd969918885, `RNS_PRIME_BITS'd390645926, `RNS_PRIME_BITS'd522676922, `RNS_PRIME_BITS'd320373698, `RNS_PRIME_BITS'd1847365274, `RNS_PRIME_BITS'd347681037, `RNS_PRIME_BITS'd1552400984, `RNS_PRIME_BITS'd596604367, `RNS_PRIME_BITS'd881136268, `RNS_PRIME_BITS'd724110489, `RNS_PRIME_BITS'd31110500, `RNS_PRIME_BITS'd1100880140, `RNS_PRIME_BITS'd1725572759, `RNS_PRIME_BITS'd425238815, `RNS_PRIME_BITS'd1857760093, `RNS_PRIME_BITS'd715601790, `RNS_PRIME_BITS'd1172573837, `RNS_PRIME_BITS'd687762618, `RNS_PRIME_BITS'd1472190862, `RNS_PRIME_BITS'd69150429, `RNS_PRIME_BITS'd100085132, `RNS_PRIME_BITS'd614244743, `RNS_PRIME_BITS'd1830179921, `RNS_PRIME_BITS'd1403519540, `RNS_PRIME_BITS'd1576410714, `RNS_PRIME_BITS'd1932282581, `RNS_PRIME_BITS'd1206867073, `RNS_PRIME_BITS'd746314798, `RNS_PRIME_BITS'd1635235279, `RNS_PRIME_BITS'd1225771145, `RNS_PRIME_BITS'd130726263, `RNS_PRIME_BITS'd372366983, `RNS_PRIME_BITS'd1064539738, `RNS_PRIME_BITS'd811256261, `RNS_PRIME_BITS'd1676468327, `RNS_PRIME_BITS'd1681719117, `RNS_PRIME_BITS'd899635798, `RNS_PRIME_BITS'd2065330097, `RNS_PRIME_BITS'd662979577, `RNS_PRIME_BITS'd1050632062, `RNS_PRIME_BITS'd794435263, `RNS_PRIME_BITS'd66648376, `RNS_PRIME_BITS'd720404290, `RNS_PRIME_BITS'd309168117, `RNS_PRIME_BITS'd1604242461, `RNS_PRIME_BITS'd1829857110, `RNS_PRIME_BITS'd982359344, `RNS_PRIME_BITS'd326449776, `RNS_PRIME_BITS'd1601120085, `RNS_PRIME_BITS'd475235749, `RNS_PRIME_BITS'd97394646, `RNS_PRIME_BITS'd991236607}
};

parameter B_BASIS_poly twist_factor_b   = '{
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd982714381, `RNS_PRIME_BITS'd1654849230, `RNS_PRIME_BITS'd478051828, `RNS_PRIME_BITS'd356657619, `RNS_PRIME_BITS'd1920663579, `RNS_PRIME_BITS'd302866737, `RNS_PRIME_BITS'd351262005, `RNS_PRIME_BITS'd532016628, `RNS_PRIME_BITS'd1151501468, `RNS_PRIME_BITS'd652946039, `RNS_PRIME_BITS'd1144091943, `RNS_PRIME_BITS'd1233595480, `RNS_PRIME_BITS'd327413943, `RNS_PRIME_BITS'd849304041, `RNS_PRIME_BITS'd385268797, `RNS_PRIME_BITS'd1929740512, `RNS_PRIME_BITS'd1437307346, `RNS_PRIME_BITS'd1054516963, `RNS_PRIME_BITS'd2052121271, `RNS_PRIME_BITS'd470080841, `RNS_PRIME_BITS'd1579045017, `RNS_PRIME_BITS'd297821259, `RNS_PRIME_BITS'd641843845, `RNS_PRIME_BITS'd99841913, `RNS_PRIME_BITS'd444118214, `RNS_PRIME_BITS'd1094401579, `RNS_PRIME_BITS'd936096522, `RNS_PRIME_BITS'd123364587, `RNS_PRIME_BITS'd456798682, `RNS_PRIME_BITS'd371148888, `RNS_PRIME_BITS'd958225700, `RNS_PRIME_BITS'd368900981, `RNS_PRIME_BITS'd906812118, `RNS_PRIME_BITS'd27942223, `RNS_PRIME_BITS'd895294767, `RNS_PRIME_BITS'd1022769805, `RNS_PRIME_BITS'd1552017062, `RNS_PRIME_BITS'd51446398, `RNS_PRIME_BITS'd199576301, `RNS_PRIME_BITS'd1898245248, `RNS_PRIME_BITS'd1467943930, `RNS_PRIME_BITS'd1732476368, `RNS_PRIME_BITS'd559257721, `RNS_PRIME_BITS'd1631487701, `RNS_PRIME_BITS'd1721817336, `RNS_PRIME_BITS'd421878258, `RNS_PRIME_BITS'd557994804, `RNS_PRIME_BITS'd304649431, `RNS_PRIME_BITS'd8907008, `RNS_PRIME_BITS'd271032415, `RNS_PRIME_BITS'd1720040104, `RNS_PRIME_BITS'd1766152386, `RNS_PRIME_BITS'd809081996, `RNS_PRIME_BITS'd1651675396, `RNS_PRIME_BITS'd1331311885, `RNS_PRIME_BITS'd769115895, `RNS_PRIME_BITS'd1990768752, `RNS_PRIME_BITS'd1644425917, `RNS_PRIME_BITS'd1206592301, `RNS_PRIME_BITS'd1688834505, `RNS_PRIME_BITS'd1022667949, `RNS_PRIME_BITS'd826531416, `RNS_PRIME_BITS'd423155928},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd561201457, `RNS_PRIME_BITS'd318222520, `RNS_PRIME_BITS'd1438809348, `RNS_PRIME_BITS'd1828267041, `RNS_PRIME_BITS'd1617885585, `RNS_PRIME_BITS'd1310190713, `RNS_PRIME_BITS'd1915188815, `RNS_PRIME_BITS'd1346436954, `RNS_PRIME_BITS'd804641710, `RNS_PRIME_BITS'd1430678598, `RNS_PRIME_BITS'd1654629824, `RNS_PRIME_BITS'd400618345, `RNS_PRIME_BITS'd1866406664, `RNS_PRIME_BITS'd5588299, `RNS_PRIME_BITS'd120346045, `RNS_PRIME_BITS'd80763692, `RNS_PRIME_BITS'd545997482, `RNS_PRIME_BITS'd983104082, `RNS_PRIME_BITS'd2097368234, `RNS_PRIME_BITS'd918812250, `RNS_PRIME_BITS'd2055579709, `RNS_PRIME_BITS'd1980041940, `RNS_PRIME_BITS'd1139003082, `RNS_PRIME_BITS'd159606694, `RNS_PRIME_BITS'd820749293, `RNS_PRIME_BITS'd1979993210, `RNS_PRIME_BITS'd2126679887, `RNS_PRIME_BITS'd229579563, `RNS_PRIME_BITS'd1169203214, `RNS_PRIME_BITS'd1458564334, `RNS_PRIME_BITS'd1357775805, `RNS_PRIME_BITS'd1776948932, `RNS_PRIME_BITS'd1955170315, `RNS_PRIME_BITS'd1966586531, `RNS_PRIME_BITS'd110672867, `RNS_PRIME_BITS'd1050480888, `RNS_PRIME_BITS'd1649403189, `RNS_PRIME_BITS'd554085691, `RNS_PRIME_BITS'd775123075, `RNS_PRIME_BITS'd1464394521, `RNS_PRIME_BITS'd1992441198, `RNS_PRIME_BITS'd1295673068, `RNS_PRIME_BITS'd1767109925, `RNS_PRIME_BITS'd1096154473, `RNS_PRIME_BITS'd767563666, `RNS_PRIME_BITS'd674822329, `RNS_PRIME_BITS'd1072848871, `RNS_PRIME_BITS'd552851043, `RNS_PRIME_BITS'd1274432900, `RNS_PRIME_BITS'd1263489667, `RNS_PRIME_BITS'd885989717, `RNS_PRIME_BITS'd236666624, `RNS_PRIME_BITS'd1923634752, `RNS_PRIME_BITS'd147052478, `RNS_PRIME_BITS'd773740556, `RNS_PRIME_BITS'd1915037, `RNS_PRIME_BITS'd1795377192, `RNS_PRIME_BITS'd674188376, `RNS_PRIME_BITS'd1038169980, `RNS_PRIME_BITS'd155056032, `RNS_PRIME_BITS'd1063723561, `RNS_PRIME_BITS'd552348229, `RNS_PRIME_BITS'd2022047502},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd2030504833, `RNS_PRIME_BITS'd458644985, `RNS_PRIME_BITS'd1933006424, `RNS_PRIME_BITS'd2042051371, `RNS_PRIME_BITS'd734171544, `RNS_PRIME_BITS'd2001209167, `RNS_PRIME_BITS'd1270889040, `RNS_PRIME_BITS'd662532888, `RNS_PRIME_BITS'd332110078, `RNS_PRIME_BITS'd586122886, `RNS_PRIME_BITS'd1868204885, `RNS_PRIME_BITS'd633289293, `RNS_PRIME_BITS'd1828476394, `RNS_PRIME_BITS'd1282347525, `RNS_PRIME_BITS'd679192186, `RNS_PRIME_BITS'd1110746654, `RNS_PRIME_BITS'd1048891790, `RNS_PRIME_BITS'd595179583, `RNS_PRIME_BITS'd1124820764, `RNS_PRIME_BITS'd1315499404, `RNS_PRIME_BITS'd674452159, `RNS_PRIME_BITS'd1801404655, `RNS_PRIME_BITS'd1493917469, `RNS_PRIME_BITS'd1314416481, `RNS_PRIME_BITS'd1952643917, `RNS_PRIME_BITS'd1368761486, `RNS_PRIME_BITS'd190758143, `RNS_PRIME_BITS'd1292695071, `RNS_PRIME_BITS'd326439411, `RNS_PRIME_BITS'd517075660, `RNS_PRIME_BITS'd611103098, `RNS_PRIME_BITS'd584149928, `RNS_PRIME_BITS'd140317819, `RNS_PRIME_BITS'd855293400, `RNS_PRIME_BITS'd714603448, `RNS_PRIME_BITS'd1486683312, `RNS_PRIME_BITS'd240212080, `RNS_PRIME_BITS'd840596094, `RNS_PRIME_BITS'd368477724, `RNS_PRIME_BITS'd732592157, `RNS_PRIME_BITS'd1047139254, `RNS_PRIME_BITS'd1079673294, `RNS_PRIME_BITS'd1351312793, `RNS_PRIME_BITS'd1594888548, `RNS_PRIME_BITS'd1273959981, `RNS_PRIME_BITS'd196565656, `RNS_PRIME_BITS'd1394641272, `RNS_PRIME_BITS'd500041537, `RNS_PRIME_BITS'd713754135, `RNS_PRIME_BITS'd1873914868, `RNS_PRIME_BITS'd1078246245, `RNS_PRIME_BITS'd514903787, `RNS_PRIME_BITS'd1737225677, `RNS_PRIME_BITS'd1438162619, `RNS_PRIME_BITS'd1755701290, `RNS_PRIME_BITS'd657916126, `RNS_PRIME_BITS'd743489674, `RNS_PRIME_BITS'd970993592, `RNS_PRIME_BITS'd1544729701, `RNS_PRIME_BITS'd677137612, `RNS_PRIME_BITS'd1980951143, `RNS_PRIME_BITS'd1474472800, `RNS_PRIME_BITS'd895771398},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd520071954, `RNS_PRIME_BITS'd1659477478, `RNS_PRIME_BITS'd380013956, `RNS_PRIME_BITS'd532048860, `RNS_PRIME_BITS'd1587022193, `RNS_PRIME_BITS'd678117384, `RNS_PRIME_BITS'd646964512, `RNS_PRIME_BITS'd1599846131, `RNS_PRIME_BITS'd492774328, `RNS_PRIME_BITS'd1813223460, `RNS_PRIME_BITS'd2035977623, `RNS_PRIME_BITS'd451198491, `RNS_PRIME_BITS'd1649721566, `RNS_PRIME_BITS'd2112063758, `RNS_PRIME_BITS'd730453618, `RNS_PRIME_BITS'd1888511225, `RNS_PRIME_BITS'd1946521804, `RNS_PRIME_BITS'd1078093079, `RNS_PRIME_BITS'd1326701425, `RNS_PRIME_BITS'd734192161, `RNS_PRIME_BITS'd1770001053, `RNS_PRIME_BITS'd1913561989, `RNS_PRIME_BITS'd965099418, `RNS_PRIME_BITS'd2125349561, `RNS_PRIME_BITS'd2020087064, `RNS_PRIME_BITS'd1790284840, `RNS_PRIME_BITS'd653091537, `RNS_PRIME_BITS'd131782201, `RNS_PRIME_BITS'd1893247609, `RNS_PRIME_BITS'd303751980, `RNS_PRIME_BITS'd1334847884, `RNS_PRIME_BITS'd873118585, `RNS_PRIME_BITS'd249386706, `RNS_PRIME_BITS'd2042384205, `RNS_PRIME_BITS'd1211271110, `RNS_PRIME_BITS'd499906752, `RNS_PRIME_BITS'd1757234669, `RNS_PRIME_BITS'd393905830, `RNS_PRIME_BITS'd1693926536, `RNS_PRIME_BITS'd780663828, `RNS_PRIME_BITS'd329767801, `RNS_PRIME_BITS'd2044280699, `RNS_PRIME_BITS'd379354092, `RNS_PRIME_BITS'd1987906920, `RNS_PRIME_BITS'd1075761591, `RNS_PRIME_BITS'd1790217672, `RNS_PRIME_BITS'd1753588508, `RNS_PRIME_BITS'd2052067642, `RNS_PRIME_BITS'd88328166, `RNS_PRIME_BITS'd102380589, `RNS_PRIME_BITS'd1561618962, `RNS_PRIME_BITS'd1443630163, `RNS_PRIME_BITS'd1636333534, `RNS_PRIME_BITS'd2056193828, `RNS_PRIME_BITS'd1878383483, `RNS_PRIME_BITS'd763768649, `RNS_PRIME_BITS'd1663859725, `RNS_PRIME_BITS'd1883950119, `RNS_PRIME_BITS'd1765983319, `RNS_PRIME_BITS'd1170752224, `RNS_PRIME_BITS'd1028658040, `RNS_PRIME_BITS'd581664342, `RNS_PRIME_BITS'd164737598},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1910348564, `RNS_PRIME_BITS'd221897449, `RNS_PRIME_BITS'd367995126, `RNS_PRIME_BITS'd1539132485, `RNS_PRIME_BITS'd2051390243, `RNS_PRIME_BITS'd2024510820, `RNS_PRIME_BITS'd1441807459, `RNS_PRIME_BITS'd2041325775, `RNS_PRIME_BITS'd101596083, `RNS_PRIME_BITS'd411860025, `RNS_PRIME_BITS'd1825753344, `RNS_PRIME_BITS'd1284434959, `RNS_PRIME_BITS'd341435820, `RNS_PRIME_BITS'd323800841, `RNS_PRIME_BITS'd959857878, `RNS_PRIME_BITS'd747078255, `RNS_PRIME_BITS'd172892730, `RNS_PRIME_BITS'd1581201429, `RNS_PRIME_BITS'd285618846, `RNS_PRIME_BITS'd498026890, `RNS_PRIME_BITS'd1516662357, `RNS_PRIME_BITS'd743336322, `RNS_PRIME_BITS'd221590400, `RNS_PRIME_BITS'd807294136, `RNS_PRIME_BITS'd1720419235, `RNS_PRIME_BITS'd2108289477, `RNS_PRIME_BITS'd1402153400, `RNS_PRIME_BITS'd1557026756, `RNS_PRIME_BITS'd486052227, `RNS_PRIME_BITS'd639432542, `RNS_PRIME_BITS'd566734447, `RNS_PRIME_BITS'd1361170515, `RNS_PRIME_BITS'd1756055478, `RNS_PRIME_BITS'd1707467875, `RNS_PRIME_BITS'd1147352387, `RNS_PRIME_BITS'd1986920445, `RNS_PRIME_BITS'd594637207, `RNS_PRIME_BITS'd1120665741, `RNS_PRIME_BITS'd914203855, `RNS_PRIME_BITS'd1967509349, `RNS_PRIME_BITS'd1977879822, `RNS_PRIME_BITS'd1932873997, `RNS_PRIME_BITS'd902553616, `RNS_PRIME_BITS'd1275904696, `RNS_PRIME_BITS'd187303824, `RNS_PRIME_BITS'd1691018214, `RNS_PRIME_BITS'd2146447664, `RNS_PRIME_BITS'd2080135103, `RNS_PRIME_BITS'd690462842, `RNS_PRIME_BITS'd466893867, `RNS_PRIME_BITS'd1038541210, `RNS_PRIME_BITS'd1022960172, `RNS_PRIME_BITS'd1108497895, `RNS_PRIME_BITS'd171133878, `RNS_PRIME_BITS'd1121975700, `RNS_PRIME_BITS'd1239138918, `RNS_PRIME_BITS'd58964999, `RNS_PRIME_BITS'd1584543981, `RNS_PRIME_BITS'd1014783106, `RNS_PRIME_BITS'd319429885, `RNS_PRIME_BITS'd77300856, `RNS_PRIME_BITS'd2100968896, `RNS_PRIME_BITS'd538728578},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1111366840, `RNS_PRIME_BITS'd1817702166, `RNS_PRIME_BITS'd308654393, `RNS_PRIME_BITS'd1902036916, `RNS_PRIME_BITS'd1514881435, `RNS_PRIME_BITS'd203341575, `RNS_PRIME_BITS'd1364034874, `RNS_PRIME_BITS'd1781417128, `RNS_PRIME_BITS'd1866997580, `RNS_PRIME_BITS'd337893308, `RNS_PRIME_BITS'd859229142, `RNS_PRIME_BITS'd181333865, `RNS_PRIME_BITS'd162479211, `RNS_PRIME_BITS'd1144062347, `RNS_PRIME_BITS'd1296633865, `RNS_PRIME_BITS'd1071833897, `RNS_PRIME_BITS'd1132496960, `RNS_PRIME_BITS'd265094956, `RNS_PRIME_BITS'd1422611, `RNS_PRIME_BITS'd536379334, `RNS_PRIME_BITS'd1941747448, `RNS_PRIME_BITS'd987777415, `RNS_PRIME_BITS'd1196073590, `RNS_PRIME_BITS'd2062390131, `RNS_PRIME_BITS'd1850634582, `RNS_PRIME_BITS'd1033810328, `RNS_PRIME_BITS'd1801237427, `RNS_PRIME_BITS'd1520994666, `RNS_PRIME_BITS'd1746039191, `RNS_PRIME_BITS'd729791605, `RNS_PRIME_BITS'd1779837071, `RNS_PRIME_BITS'd1162711167, `RNS_PRIME_BITS'd915333332, `RNS_PRIME_BITS'd1299152479, `RNS_PRIME_BITS'd1301194870, `RNS_PRIME_BITS'd1980475697, `RNS_PRIME_BITS'd988918344, `RNS_PRIME_BITS'd881125819, `RNS_PRIME_BITS'd237869749, `RNS_PRIME_BITS'd1814328256, `RNS_PRIME_BITS'd627285491, `RNS_PRIME_BITS'd718059950, `RNS_PRIME_BITS'd1567408049, `RNS_PRIME_BITS'd45733247, `RNS_PRIME_BITS'd1822384920, `RNS_PRIME_BITS'd1758326586, `RNS_PRIME_BITS'd1454548222, `RNS_PRIME_BITS'd1467683836, `RNS_PRIME_BITS'd630505524, `RNS_PRIME_BITS'd275250926, `RNS_PRIME_BITS'd770159278, `RNS_PRIME_BITS'd1343151649, `RNS_PRIME_BITS'd136842044, `RNS_PRIME_BITS'd103088552, `RNS_PRIME_BITS'd898174659, `RNS_PRIME_BITS'd218696274, `RNS_PRIME_BITS'd1758502347, `RNS_PRIME_BITS'd194569702, `RNS_PRIME_BITS'd1833115473, `RNS_PRIME_BITS'd2146875856, `RNS_PRIME_BITS'd1385487051, `RNS_PRIME_BITS'd594047528, `RNS_PRIME_BITS'd91096341},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1316470784, `RNS_PRIME_BITS'd1453892451, `RNS_PRIME_BITS'd1313726466, `RNS_PRIME_BITS'd1435226373, `RNS_PRIME_BITS'd789663591, `RNS_PRIME_BITS'd1428696568, `RNS_PRIME_BITS'd1692753891, `RNS_PRIME_BITS'd1222739369, `RNS_PRIME_BITS'd1601511596, `RNS_PRIME_BITS'd1424810859, `RNS_PRIME_BITS'd1150701755, `RNS_PRIME_BITS'd1443308359, `RNS_PRIME_BITS'd214516484, `RNS_PRIME_BITS'd908740576, `RNS_PRIME_BITS'd918632540, `RNS_PRIME_BITS'd1181774526, `RNS_PRIME_BITS'd95042921, `RNS_PRIME_BITS'd162700068, `RNS_PRIME_BITS'd922037797, `RNS_PRIME_BITS'd608940391, `RNS_PRIME_BITS'd1162784154, `RNS_PRIME_BITS'd385218143, `RNS_PRIME_BITS'd789327398, `RNS_PRIME_BITS'd1394307591, `RNS_PRIME_BITS'd541471192, `RNS_PRIME_BITS'd385488776, `RNS_PRIME_BITS'd871114005, `RNS_PRIME_BITS'd1975029035, `RNS_PRIME_BITS'd953927283, `RNS_PRIME_BITS'd220568782, `RNS_PRIME_BITS'd1814090713, `RNS_PRIME_BITS'd2018759315, `RNS_PRIME_BITS'd1392338561, `RNS_PRIME_BITS'd1860847603, `RNS_PRIME_BITS'd987706370, `RNS_PRIME_BITS'd587044175, `RNS_PRIME_BITS'd99971581, `RNS_PRIME_BITS'd649424080, `RNS_PRIME_BITS'd815239180, `RNS_PRIME_BITS'd216334037, `RNS_PRIME_BITS'd1040898177, `RNS_PRIME_BITS'd1226695548, `RNS_PRIME_BITS'd2004174612, `RNS_PRIME_BITS'd2109392002, `RNS_PRIME_BITS'd133379464, `RNS_PRIME_BITS'd1733682231, `RNS_PRIME_BITS'd2118490453, `RNS_PRIME_BITS'd353404950, `RNS_PRIME_BITS'd286276109, `RNS_PRIME_BITS'd86404339, `RNS_PRIME_BITS'd1246377055, `RNS_PRIME_BITS'd972264218, `RNS_PRIME_BITS'd350723734, `RNS_PRIME_BITS'd611788180, `RNS_PRIME_BITS'd2046419506, `RNS_PRIME_BITS'd211766403, `RNS_PRIME_BITS'd1172996175, `RNS_PRIME_BITS'd1142519638, `RNS_PRIME_BITS'd93701488, `RNS_PRIME_BITS'd1943881058, `RNS_PRIME_BITS'd1817397096, `RNS_PRIME_BITS'd752878080, `RNS_PRIME_BITS'd1545542847},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd2130228297, `RNS_PRIME_BITS'd1033346514, `RNS_PRIME_BITS'd581750232, `RNS_PRIME_BITS'd1625142860, `RNS_PRIME_BITS'd486721859, `RNS_PRIME_BITS'd571204460, `RNS_PRIME_BITS'd981144746, `RNS_PRIME_BITS'd574229214, `RNS_PRIME_BITS'd1089218493, `RNS_PRIME_BITS'd26513139, `RNS_PRIME_BITS'd2010605865, `RNS_PRIME_BITS'd341692242, `RNS_PRIME_BITS'd1506386962, `RNS_PRIME_BITS'd1816898220, `RNS_PRIME_BITS'd313660301, `RNS_PRIME_BITS'd1944313893, `RNS_PRIME_BITS'd1484566497, `RNS_PRIME_BITS'd1541045115, `RNS_PRIME_BITS'd630923484, `RNS_PRIME_BITS'd2064395269, `RNS_PRIME_BITS'd1090276043, `RNS_PRIME_BITS'd2012553244, `RNS_PRIME_BITS'd1510469846, `RNS_PRIME_BITS'd337677835, `RNS_PRIME_BITS'd1602631169, `RNS_PRIME_BITS'd972301580, `RNS_PRIME_BITS'd1727682728, `RNS_PRIME_BITS'd1168805901, `RNS_PRIME_BITS'd1956709734, `RNS_PRIME_BITS'd73418631, `RNS_PRIME_BITS'd1880750118, `RNS_PRIME_BITS'd2098452362, `RNS_PRIME_BITS'd554672634, `RNS_PRIME_BITS'd1726140753, `RNS_PRIME_BITS'd54660901, `RNS_PRIME_BITS'd818416481, `RNS_PRIME_BITS'd1747488468, `RNS_PRIME_BITS'd1455471245, `RNS_PRIME_BITS'd692845039, `RNS_PRIME_BITS'd551036518, `RNS_PRIME_BITS'd1927967098, `RNS_PRIME_BITS'd319374927, `RNS_PRIME_BITS'd1915883062, `RNS_PRIME_BITS'd1049625500, `RNS_PRIME_BITS'd184438272, `RNS_PRIME_BITS'd1734877556, `RNS_PRIME_BITS'd1685711725, `RNS_PRIME_BITS'd1945521432, `RNS_PRIME_BITS'd1094799911, `RNS_PRIME_BITS'd353031189, `RNS_PRIME_BITS'd1813434134, `RNS_PRIME_BITS'd1923012750, `RNS_PRIME_BITS'd1158896720, `RNS_PRIME_BITS'd1273570555, `RNS_PRIME_BITS'd130023201, `RNS_PRIME_BITS'd1362281852, `RNS_PRIME_BITS'd96243187, `RNS_PRIME_BITS'd1736961913, `RNS_PRIME_BITS'd1821585998, `RNS_PRIME_BITS'd695913565, `RNS_PRIME_BITS'd694079929, `RNS_PRIME_BITS'd295372288, `RNS_PRIME_BITS'd592953865},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd1972786723, `RNS_PRIME_BITS'd1445995283, `RNS_PRIME_BITS'd1987253116, `RNS_PRIME_BITS'd501746762, `RNS_PRIME_BITS'd463114787, `RNS_PRIME_BITS'd108107719, `RNS_PRIME_BITS'd1680185572, `RNS_PRIME_BITS'd1267807369, `RNS_PRIME_BITS'd1018407763, `RNS_PRIME_BITS'd1846795101, `RNS_PRIME_BITS'd1267530456, `RNS_PRIME_BITS'd246731728, `RNS_PRIME_BITS'd1125681298, `RNS_PRIME_BITS'd1797675798, `RNS_PRIME_BITS'd1117135201, `RNS_PRIME_BITS'd849564324, `RNS_PRIME_BITS'd1508207091, `RNS_PRIME_BITS'd251058699, `RNS_PRIME_BITS'd1729285507, `RNS_PRIME_BITS'd796429192, `RNS_PRIME_BITS'd2067686905, `RNS_PRIME_BITS'd1979833503, `RNS_PRIME_BITS'd270694143, `RNS_PRIME_BITS'd132886023, `RNS_PRIME_BITS'd1160547813, `RNS_PRIME_BITS'd464279201, `RNS_PRIME_BITS'd1152260240, `RNS_PRIME_BITS'd422202768, `RNS_PRIME_BITS'd48756347, `RNS_PRIME_BITS'd1842850055, `RNS_PRIME_BITS'd583666609, `RNS_PRIME_BITS'd1282120144, `RNS_PRIME_BITS'd1803248469, `RNS_PRIME_BITS'd327226555, `RNS_PRIME_BITS'd819125480, `RNS_PRIME_BITS'd35025808, `RNS_PRIME_BITS'd1882163270, `RNS_PRIME_BITS'd458116540, `RNS_PRIME_BITS'd768852906, `RNS_PRIME_BITS'd1945334986, `RNS_PRIME_BITS'd1632011555, `RNS_PRIME_BITS'd1006104391, `RNS_PRIME_BITS'd1568208839, `RNS_PRIME_BITS'd1719836841, `RNS_PRIME_BITS'd1461368271, `RNS_PRIME_BITS'd416072182, `RNS_PRIME_BITS'd726102973, `RNS_PRIME_BITS'd1970029940, `RNS_PRIME_BITS'd1229835195, `RNS_PRIME_BITS'd611355256, `RNS_PRIME_BITS'd792897446, `RNS_PRIME_BITS'd108303762, `RNS_PRIME_BITS'd928987687, `RNS_PRIME_BITS'd2141801975, `RNS_PRIME_BITS'd1602925057, `RNS_PRIME_BITS'd1719197983, `RNS_PRIME_BITS'd1842468980, `RNS_PRIME_BITS'd335514896, `RNS_PRIME_BITS'd1974242872, `RNS_PRIME_BITS'd1405654688, `RNS_PRIME_BITS'd1947249161, `RNS_PRIME_BITS'd862305235, `RNS_PRIME_BITS'd516818747},
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd601347331, `RNS_PRIME_BITS'd330138710, `RNS_PRIME_BITS'd1006948292, `RNS_PRIME_BITS'd211376156, `RNS_PRIME_BITS'd15801270, `RNS_PRIME_BITS'd97888807, `RNS_PRIME_BITS'd1297233476, `RNS_PRIME_BITS'd125361803, `RNS_PRIME_BITS'd1327782020, `RNS_PRIME_BITS'd774401595, `RNS_PRIME_BITS'd993630259, `RNS_PRIME_BITS'd830621476, `RNS_PRIME_BITS'd213719977, `RNS_PRIME_BITS'd1784673181, `RNS_PRIME_BITS'd244734214, `RNS_PRIME_BITS'd634071871, `RNS_PRIME_BITS'd1357050316, `RNS_PRIME_BITS'd850930788, `RNS_PRIME_BITS'd1908735073, `RNS_PRIME_BITS'd855303704, `RNS_PRIME_BITS'd892337725, `RNS_PRIME_BITS'd518922129, `RNS_PRIME_BITS'd120244624, `RNS_PRIME_BITS'd590119148, `RNS_PRIME_BITS'd1858954969, `RNS_PRIME_BITS'd627138487, `RNS_PRIME_BITS'd886133038, `RNS_PRIME_BITS'd44695371, `RNS_PRIME_BITS'd747272326, `RNS_PRIME_BITS'd1029685765, `RNS_PRIME_BITS'd1598964437, `RNS_PRIME_BITS'd764279395, `RNS_PRIME_BITS'd973858991, `RNS_PRIME_BITS'd1314367513, `RNS_PRIME_BITS'd1786870076, `RNS_PRIME_BITS'd996800473, `RNS_PRIME_BITS'd456097637, `RNS_PRIME_BITS'd1687641260, `RNS_PRIME_BITS'd460818202, `RNS_PRIME_BITS'd1264514118, `RNS_PRIME_BITS'd1401930789, `RNS_PRIME_BITS'd703232155, `RNS_PRIME_BITS'd799915249, `RNS_PRIME_BITS'd279176347, `RNS_PRIME_BITS'd313264892, `RNS_PRIME_BITS'd1441277666, `RNS_PRIME_BITS'd223845845, `RNS_PRIME_BITS'd2061554458, `RNS_PRIME_BITS'd1665960726, `RNS_PRIME_BITS'd990739525, `RNS_PRIME_BITS'd76817238, `RNS_PRIME_BITS'd616062626, `RNS_PRIME_BITS'd1278419481, `RNS_PRIME_BITS'd1138746994, `RNS_PRIME_BITS'd740347681, `RNS_PRIME_BITS'd794875457, `RNS_PRIME_BITS'd1779277119, `RNS_PRIME_BITS'd1006865747, `RNS_PRIME_BITS'd1512458516, `RNS_PRIME_BITS'd520640850, `RNS_PRIME_BITS'd629079252, `RNS_PRIME_BITS'd1708924581, `RNS_PRIME_BITS'd1490950549}
};
parameter B_BASIS_poly untwist_factor_b = '{
    '{`RNS_PRIME_BITS'd2113938037, `RNS_PRIME_BITS'd798697917, `RNS_PRIME_BITS'd792395175, `RNS_PRIME_BITS'd1493976554, `RNS_PRIME_BITS'd275603109, `RNS_PRIME_BITS'd1491102736, `RNS_PRIME_BITS'd2021134738, `RNS_PRIME_BITS'd1579513695, `RNS_PRIME_BITS'd1833484025, `RNS_PRIME_BITS'd415407688, `RNS_PRIME_BITS'd108410860, `RNS_PRIME_BITS'd390012958, `RNS_PRIME_BITS'd39513013, `RNS_PRIME_BITS'd1315307254, `RNS_PRIME_BITS'd1035956851, `RNS_PRIME_BITS'd2147353437, `RNS_PRIME_BITS'd766995009, `RNS_PRIME_BITS'd1736119076, `RNS_PRIME_BITS'd1671136753, `RNS_PRIME_BITS'd1852152637, `RNS_PRIME_BITS'd679154017, `RNS_PRIME_BITS'd1903872203, `RNS_PRIME_BITS'd509803209, `RNS_PRIME_BITS'd1923228553, `RNS_PRIME_BITS'd2117832527, `RNS_PRIME_BITS'd1506837361, `RNS_PRIME_BITS'd2079579615, `RNS_PRIME_BITS'd1250823470, `RNS_PRIME_BITS'd420228658, `RNS_PRIME_BITS'd1563075904, `RNS_PRIME_BITS'd502881983, `RNS_PRIME_BITS'd724031645, `RNS_PRIME_BITS'd1772628239, `RNS_PRIME_BITS'd1192992316, `RNS_PRIME_BITS'd799510527, `RNS_PRIME_BITS'd865281393, `RNS_PRIME_BITS'd1440919025, `RNS_PRIME_BITS'd320919212, `RNS_PRIME_BITS'd1425746572, `RNS_PRIME_BITS'd194388085, `RNS_PRIME_BITS'd1911050575, `RNS_PRIME_BITS'd157744050, `RNS_PRIME_BITS'd364446835, `RNS_PRIME_BITS'd814191722, `RNS_PRIME_BITS'd294646135, `RNS_PRIME_BITS'd1813437066, `RNS_PRIME_BITS'd1157933193, `RNS_PRIME_BITS'd581524369, `RNS_PRIME_BITS'd1043594109, `RNS_PRIME_BITS'd2040809068, `RNS_PRIME_BITS'd1362467077, `RNS_PRIME_BITS'd1840385618, `RNS_PRIME_BITS'd786034799, `RNS_PRIME_BITS'd1290751872, `RNS_PRIME_BITS'd1835299179, `RNS_PRIME_BITS'd921535806, `RNS_PRIME_BITS'd1736524985, `RNS_PRIME_BITS'd1772903848, `RNS_PRIME_BITS'd1639441736, `RNS_PRIME_BITS'd875963076, `RNS_PRIME_BITS'd631964093, `RNS_PRIME_BITS'd1737368185, `RNS_PRIME_BITS'd443906989, `RNS_PRIME_BITS'd420854524},
    '{`RNS_PRIME_BITS'd2113939297, `RNS_PRIME_BITS'd438169796, `RNS_PRIME_BITS'd159142519, `RNS_PRIME_BITS'd1359117592, `RNS_PRIME_BITS'd1071324194, `RNS_PRIME_BITS'd1997054115, `RNS_PRIME_BITS'd794776015, `RNS_PRIME_BITS'd1314130912, `RNS_PRIME_BITS'd973053246, `RNS_PRIME_BITS'd390565408, `RNS_PRIME_BITS'd2078087010, `RNS_PRIME_BITS'd2117437096, `RNS_PRIME_BITS'd2143795973, `RNS_PRIME_BITS'd690802843, `RNS_PRIME_BITS'd80921750, `RNS_PRIME_BITS'd114305354, `RNS_PRIME_BITS'd1165772423, `RNS_PRIME_BITS'd1291865825, `RNS_PRIME_BITS'd1902067646, `RNS_PRIME_BITS'd591989474, `RNS_PRIME_BITS'd1358610859, `RNS_PRIME_BITS'd1213908812, `RNS_PRIME_BITS'd1456157157, `RNS_PRIME_BITS'd1512379339, `RNS_PRIME_BITS'd815983636, `RNS_PRIME_BITS'd88552478, `RNS_PRIME_BITS'd1971063340, `RNS_PRIME_BITS'd1752621452, `RNS_PRIME_BITS'd1862643389, `RNS_PRIME_BITS'd1172681457, `RNS_PRIME_BITS'd1143682806, `RNS_PRIME_BITS'd338550976, `RNS_PRIME_BITS'd106453541, `RNS_PRIME_BITS'd2025614866, `RNS_PRIME_BITS'd1520721165, `RNS_PRIME_BITS'd451495488, `RNS_PRIME_BITS'd1439260276, `RNS_PRIME_BITS'd470089507, `RNS_PRIME_BITS'd1915228943, `RNS_PRIME_BITS'd1497132433, `RNS_PRIME_BITS'd1272580642, `RNS_PRIME_BITS'd317748997, `RNS_PRIME_BITS'd640153685, `RNS_PRIME_BITS'd2014711680, `RNS_PRIME_BITS'd858062951, `RNS_PRIME_BITS'd1376521486, `RNS_PRIME_BITS'd588621655, `RNS_PRIME_BITS'd1400761654, `RNS_PRIME_BITS'd1475140116, `RNS_PRIME_BITS'd2044949706, `RNS_PRIME_BITS'd369013195, `RNS_PRIME_BITS'd239274132, `RNS_PRIME_BITS'd1369478611, `RNS_PRIME_BITS'd2121640298, `RNS_PRIME_BITS'd178973199, `RNS_PRIME_BITS'd1530938706, `RNS_PRIME_BITS'd851381315, `RNS_PRIME_BITS'd473394055, `RNS_PRIME_BITS'd1892140015, `RNS_PRIME_BITS'd545148602, `RNS_PRIME_BITS'd1078734864, `RNS_PRIME_BITS'd111736972, `RNS_PRIME_BITS'd1874084926, `RNS_PRIME_BITS'd1635406236},
    '{`RNS_PRIME_BITS'd2113939675, `RNS_PRIME_BITS'd187331160, `RNS_PRIME_BITS'd1050708499, `RNS_PRIME_BITS'd1277676961, `RNS_PRIME_BITS'd392074901, `RNS_PRIME_BITS'd1217383725, `RNS_PRIME_BITS'd1863885714, `RNS_PRIME_BITS'd323928954, `RNS_PRIME_BITS'd996358001, `RNS_PRIME_BITS'd1381860284, `RNS_PRIME_BITS'd1957249992, `RNS_PRIME_BITS'd409065623, `RNS_PRIME_BITS'd1434802343, `RNS_PRIME_BITS'd1224672529, `RNS_PRIME_BITS'd1715559177, `RNS_PRIME_BITS'd760603346, `RNS_PRIME_BITS'd25741449, `RNS_PRIME_BITS'd1857266219, `RNS_PRIME_BITS'd802239014, `RNS_PRIME_BITS'd1490051286, `RNS_PRIME_BITS'd1183045395, `RNS_PRIME_BITS'd817750688, `RNS_PRIME_BITS'd452894477, `RNS_PRIME_BITS'd1795586742, `RNS_PRIME_BITS'd961636590, `RNS_PRIME_BITS'd933771280, `RNS_PRIME_BITS'd2067250763, `RNS_PRIME_BITS'd1606867391, `RNS_PRIME_BITS'd1587391278, `RNS_PRIME_BITS'd1867891810, `RNS_PRIME_BITS'd791946393, `RNS_PRIME_BITS'd1977528817, `RNS_PRIME_BITS'd1333056578, `RNS_PRIME_BITS'd1936618199, `RNS_PRIME_BITS'd394575869, `RNS_PRIME_BITS'd1706183883, `RNS_PRIME_BITS'd1019994178, `RNS_PRIME_BITS'd2110959079, `RNS_PRIME_BITS'd448377474, `RNS_PRIME_BITS'd405699713, `RNS_PRIME_BITS'd1086763977, `RNS_PRIME_BITS'd949740882, `RNS_PRIME_BITS'd1548919159, `RNS_PRIME_BITS'd2103401360, `RNS_PRIME_BITS'd382100498, `RNS_PRIME_BITS'd921953420, `RNS_PRIME_BITS'd2104639994, `RNS_PRIME_BITS'd453375438, `RNS_PRIME_BITS'd989282524, `RNS_PRIME_BITS'd1935554307, `RNS_PRIME_BITS'd147736310, `RNS_PRIME_BITS'd1380723173, `RNS_PRIME_BITS'd426314629, `RNS_PRIME_BITS'd675455857, `RNS_PRIME_BITS'd192169418, `RNS_PRIME_BITS'd2075195857, `RNS_PRIME_BITS'd794958276, `RNS_PRIME_BITS'd517015927, `RNS_PRIME_BITS'd472050077, `RNS_PRIME_BITS'd793838922, `RNS_PRIME_BITS'd1410940662, `RNS_PRIME_BITS'd775107127, `RNS_PRIME_BITS'd1905445759, `RNS_PRIME_BITS'd1827960},
    '{`RNS_PRIME_BITS'd2113939927, `RNS_PRIME_BITS'd2077811300, `RNS_PRIME_BITS'd729112739, `RNS_PRIME_BITS'd1862984931, `RNS_PRIME_BITS'd1055454261, `RNS_PRIME_BITS'd744162357, `RNS_PRIME_BITS'd1279192758, `RNS_PRIME_BITS'd410212018, `RNS_PRIME_BITS'd290057533, `RNS_PRIME_BITS'd1950371777, `RNS_PRIME_BITS'd1175837644, `RNS_PRIME_BITS'd981070349, `RNS_PRIME_BITS'd614980717, `RNS_PRIME_BITS'd579582540, `RNS_PRIME_BITS'd1508357394, `RNS_PRIME_BITS'd1273694749, `RNS_PRIME_BITS'd1914103360, `RNS_PRIME_BITS'd912129036, `RNS_PRIME_BITS'd240464665, `RNS_PRIME_BITS'd1828694336, `RNS_PRIME_BITS'd1311123035, `RNS_PRIME_BITS'd1470475081, `RNS_PRIME_BITS'd1947779633, `RNS_PRIME_BITS'd1907459693, `RNS_PRIME_BITS'd658894168, `RNS_PRIME_BITS'd241969214, `RNS_PRIME_BITS'd1268920098, `RNS_PRIME_BITS'd1482500299, `RNS_PRIME_BITS'd2139683486, `RNS_PRIME_BITS'd182401501, `RNS_PRIME_BITS'd404297573, `RNS_PRIME_BITS'd600086169, `RNS_PRIME_BITS'd1898969837, `RNS_PRIME_BITS'd381798226, `RNS_PRIME_BITS'd1471656364, `RNS_PRIME_BITS'd1883030321, `RNS_PRIME_BITS'd1910553218, `RNS_PRIME_BITS'd560223679, `RNS_PRIME_BITS'd1314210880, `RNS_PRIME_BITS'd773746588, `RNS_PRIME_BITS'd1879403728, `RNS_PRIME_BITS'd857339974, `RNS_PRIME_BITS'd137873604, `RNS_PRIME_BITS'd945427192, `RNS_PRIME_BITS'd1095830114, `RNS_PRIME_BITS'd1623445789, `RNS_PRIME_BITS'd754910642, `RNS_PRIME_BITS'd372240821, `RNS_PRIME_BITS'd1883104327, `RNS_PRIME_BITS'd1666316763, `RNS_PRIME_BITS'd436763432, `RNS_PRIME_BITS'd980861161, `RNS_PRIME_BITS'd898924278, `RNS_PRIME_BITS'd739943696, `RNS_PRIME_BITS'd1179634056, `RNS_PRIME_BITS'd1871358114, `RNS_PRIME_BITS'd1686287107, `RNS_PRIME_BITS'd1063638444, `RNS_PRIME_BITS'd257841232, `RNS_PRIME_BITS'd1619378277, `RNS_PRIME_BITS'd931215593, `RNS_PRIME_BITS'd128280690, `RNS_PRIME_BITS'd1249145541, `RNS_PRIME_BITS'd595856712},
    '{`RNS_PRIME_BITS'd2113940305, `RNS_PRIME_BITS'd58691582, `RNS_PRIME_BITS'd2114667274, `RNS_PRIME_BITS'd1877850223, `RNS_PRIME_BITS'd2041839997, `RNS_PRIME_BITS'd51253230, `RNS_PRIME_BITS'd1485198861, `RNS_PRIME_BITS'd233960928, `RNS_PRIME_BITS'd1255713559, `RNS_PRIME_BITS'd653561290, `RNS_PRIME_BITS'd1809274866, `RNS_PRIME_BITS'd1291309433, `RNS_PRIME_BITS'd1460419000, `RNS_PRIME_BITS'd856192602, `RNS_PRIME_BITS'd1435552928, `RNS_PRIME_BITS'd1935378783, `RNS_PRIME_BITS'd2081438194, `RNS_PRIME_BITS'd1577082940, `RNS_PRIME_BITS'd1248652945, `RNS_PRIME_BITS'd533947106, `RNS_PRIME_BITS'd1859122038, `RNS_PRIME_BITS'd522771328, `RNS_PRIME_BITS'd406008748, `RNS_PRIME_BITS'd438860140, `RNS_PRIME_BITS'd1210778163, `RNS_PRIME_BITS'd489034685, `RNS_PRIME_BITS'd418699502, `RNS_PRIME_BITS'd762464778, `RNS_PRIME_BITS'd2015785457, `RNS_PRIME_BITS'd82736443, `RNS_PRIME_BITS'd1147732095, `RNS_PRIME_BITS'd1784510466, `RNS_PRIME_BITS'd616269263, `RNS_PRIME_BITS'd1568211351, `RNS_PRIME_BITS'd996647107, `RNS_PRIME_BITS'd93069258, `RNS_PRIME_BITS'd109889889, `RNS_PRIME_BITS'd1857149402, `RNS_PRIME_BITS'd134831017, `RNS_PRIME_BITS'd1147529730, `RNS_PRIME_BITS'd1866444078, `RNS_PRIME_BITS'd2144032563, `RNS_PRIME_BITS'd55494586, `RNS_PRIME_BITS'd680948919, `RNS_PRIME_BITS'd327764410, `RNS_PRIME_BITS'd1002175446, `RNS_PRIME_BITS'd679940496, `RNS_PRIME_BITS'd1943465816, `RNS_PRIME_BITS'd1565393479, `RNS_PRIME_BITS'd723203597, `RNS_PRIME_BITS'd296932084, `RNS_PRIME_BITS'd1471067818, `RNS_PRIME_BITS'd483249824, `RNS_PRIME_BITS'd2118967517, `RNS_PRIME_BITS'd1906177344, `RNS_PRIME_BITS'd1709697570, `RNS_PRIME_BITS'd471423405, `RNS_PRIME_BITS'd1151883039, `RNS_PRIME_BITS'd1176332907, `RNS_PRIME_BITS'd1142358308, `RNS_PRIME_BITS'd143724095, `RNS_PRIME_BITS'd1806198909, `RNS_PRIME_BITS'd1372271781, `RNS_PRIME_BITS'd641242964},
    '{`RNS_PRIME_BITS'd2113941061, `RNS_PRIME_BITS'd703223640, `RNS_PRIME_BITS'd1332902808, `RNS_PRIME_BITS'd347452585, `RNS_PRIME_BITS'd503328985, `RNS_PRIME_BITS'd541786111, `RNS_PRIME_BITS'd1272035409, `RNS_PRIME_BITS'd341624221, `RNS_PRIME_BITS'd600566031, `RNS_PRIME_BITS'd86629881, `RNS_PRIME_BITS'd1340574042, `RNS_PRIME_BITS'd2011139044, `RNS_PRIME_BITS'd1086315716, `RNS_PRIME_BITS'd1531478782, `RNS_PRIME_BITS'd1539211725, `RNS_PRIME_BITS'd1734988592, `RNS_PRIME_BITS'd1990344641, `RNS_PRIME_BITS'd2057659125, `RNS_PRIME_BITS'd1918694108, `RNS_PRIME_BITS'd776836116, `RNS_PRIME_BITS'd2113226479, `RNS_PRIME_BITS'd1619685630, `RNS_PRIME_BITS'd1532292834, `RNS_PRIME_BITS'd1701484285, `RNS_PRIME_BITS'd2119146802, `RNS_PRIME_BITS'd1774678146, `RNS_PRIME_BITS'd1965954990, `RNS_PRIME_BITS'd252985111, `RNS_PRIME_BITS'd1613231448, `RNS_PRIME_BITS'd1791618311, `RNS_PRIME_BITS'd1019893963, `RNS_PRIME_BITS'd656790317, `RNS_PRIME_BITS'd2095773699, `RNS_PRIME_BITS'd475509346, `RNS_PRIME_BITS'd1766991867, `RNS_PRIME_BITS'd744474398, `RNS_PRIME_BITS'd1385528499, `RNS_PRIME_BITS'd1683141286, `RNS_PRIME_BITS'd789157594, `RNS_PRIME_BITS'd709285475, `RNS_PRIME_BITS'd1679060775, `RNS_PRIME_BITS'd1793260831, `RNS_PRIME_BITS'd219448318, `RNS_PRIME_BITS'd1848718917, `RNS_PRIME_BITS'd192946793, `RNS_PRIME_BITS'd637515552, `RNS_PRIME_BITS'd1472261172, `RNS_PRIME_BITS'd2129800416, `RNS_PRIME_BITS'd1358992016, `RNS_PRIME_BITS'd281731676, `RNS_PRIME_BITS'd351224846, `RNS_PRIME_BITS'd1440309923, `RNS_PRIME_BITS'd1372906079, `RNS_PRIME_BITS'd724776185, `RNS_PRIME_BITS'd2007997618, `RNS_PRIME_BITS'd373483603, `RNS_PRIME_BITS'd1314350158, `RNS_PRIME_BITS'd1924854916, `RNS_PRIME_BITS'd231705128, `RNS_PRIME_BITS'd882304718, `RNS_PRIME_BITS'd1715120914, `RNS_PRIME_BITS'd1907790616, `RNS_PRIME_BITS'd709800044, `RNS_PRIME_BITS'd1861693614},
    '{`RNS_PRIME_BITS'd2113941565, `RNS_PRIME_BITS'd2089792458, `RNS_PRIME_BITS'd2135732473, `RNS_PRIME_BITS'd1313788291, `RNS_PRIME_BITS'd1110484211, `RNS_PRIME_BITS'd1609158059, `RNS_PRIME_BITS'd720349947, `RNS_PRIME_BITS'd484991355, `RNS_PRIME_BITS'd97355034, `RNS_PRIME_BITS'd1645756096, `RNS_PRIME_BITS'd661533370, `RNS_PRIME_BITS'd732721758, `RNS_PRIME_BITS'd857228700, `RNS_PRIME_BITS'd1020718827, `RNS_PRIME_BITS'd1709935961, `RNS_PRIME_BITS'd431737100, `RNS_PRIME_BITS'd732679864, `RNS_PRIME_BITS'd671545775, `RNS_PRIME_BITS'd1818415756, `RNS_PRIME_BITS'd266352970, `RNS_PRIME_BITS'd34150006, `RNS_PRIME_BITS'd639777332, `RNS_PRIME_BITS'd1994110563, `RNS_PRIME_BITS'd17290594, `RNS_PRIME_BITS'd701266969, `RNS_PRIME_BITS'd389917424, `RNS_PRIME_BITS'd526726797, `RNS_PRIME_BITS'd2045270253, `RNS_PRIME_BITS'd494146855, `RNS_PRIME_BITS'd51676344, `RNS_PRIME_BITS'd1682210285, `RNS_PRIME_BITS'd11799338, `RNS_PRIME_BITS'd605994818, `RNS_PRIME_BITS'd810520533, `RNS_PRIME_BITS'd466318405, `RNS_PRIME_BITS'd1696380915, `RNS_PRIME_BITS'd1411989176, `RNS_PRIME_BITS'd691036032, `RNS_PRIME_BITS'd262413762, `RNS_PRIME_BITS'd796850585, `RNS_PRIME_BITS'd213096340, `RNS_PRIME_BITS'd1262742624, `RNS_PRIME_BITS'd1034174435, `RNS_PRIME_BITS'd854251826, `RNS_PRIME_BITS'd1299115799, `RNS_PRIME_BITS'd1227114396, `RNS_PRIME_BITS'd1205424420, `RNS_PRIME_BITS'd1374254703, `RNS_PRIME_BITS'd2061921710, `RNS_PRIME_BITS'd925175951, `RNS_PRIME_BITS'd1059549025, `RNS_PRIME_BITS'd130866692, `RNS_PRIME_BITS'd212330703, `RNS_PRIME_BITS'd1961743338, `RNS_PRIME_BITS'd1420586335, `RNS_PRIME_BITS'd1451380014, `RNS_PRIME_BITS'd1356634446, `RNS_PRIME_BITS'd1147962701, `RNS_PRIME_BITS'd1856735785, `RNS_PRIME_BITS'd1296291999, `RNS_PRIME_BITS'd145347728, `RNS_PRIME_BITS'd46582280, `RNS_PRIME_BITS'd1151694911, `RNS_PRIME_BITS'd2126926337},
    '{`RNS_PRIME_BITS'd2113942321, `RNS_PRIME_BITS'd292726856, `RNS_PRIME_BITS'd2142881769, `RNS_PRIME_BITS'd1901769482, `RNS_PRIME_BITS'd962210911, `RNS_PRIME_BITS'd441302679, `RNS_PRIME_BITS'd1885474451, `RNS_PRIME_BITS'd1709782841, `RNS_PRIME_BITS'd1991992747, `RNS_PRIME_BITS'd1105271508, `RNS_PRIME_BITS'd1959824221, `RNS_PRIME_BITS'd518766479, `RNS_PRIME_BITS'd439717886, `RNS_PRIME_BITS'd709867172, `RNS_PRIME_BITS'd699131328, `RNS_PRIME_BITS'd1291524712, `RNS_PRIME_BITS'd774912588, `RNS_PRIME_BITS'd1483619555, `RNS_PRIME_BITS'd1717733819, `RNS_PRIME_BITS'd2144615113, `RNS_PRIME_BITS'd923129522, `RNS_PRIME_BITS'd1782014888, `RNS_PRIME_BITS'd498329367, `RNS_PRIME_BITS'd1916044635, `RNS_PRIME_BITS'd1266466375, `RNS_PRIME_BITS'd1566242377, `RNS_PRIME_BITS'd413468582, `RNS_PRIME_BITS'd643788293, `RNS_PRIME_BITS'd1094515363, `RNS_PRIME_BITS'd1240667604, `RNS_PRIME_BITS'd543457931, `RNS_PRIME_BITS'd1937502361, `RNS_PRIME_BITS'd302758082, `RNS_PRIME_BITS'd1245689600, `RNS_PRIME_BITS'd233735314, `RNS_PRIME_BITS'd1244502731, `RNS_PRIME_BITS'd417947728, `RNS_PRIME_BITS'd1315190558, `RNS_PRIME_BITS'd387463468, `RNS_PRIME_BITS'd8513528, `RNS_PRIME_BITS'd363824824, `RNS_PRIME_BITS'd714600989, `RNS_PRIME_BITS'd908083776, `RNS_PRIME_BITS'd352065477, `RNS_PRIME_BITS'd135517024, `RNS_PRIME_BITS'd929671741, `RNS_PRIME_BITS'd1955644931, `RNS_PRIME_BITS'd1084106769, `RNS_PRIME_BITS'd1211141776, `RNS_PRIME_BITS'd431309378, `RNS_PRIME_BITS'd1448015126, `RNS_PRIME_BITS'd580446224, `RNS_PRIME_BITS'd598644579, `RNS_PRIME_BITS'd1344324524, `RNS_PRIME_BITS'd1710872373, `RNS_PRIME_BITS'd2029814002, `RNS_PRIME_BITS'd997666869, `RNS_PRIME_BITS'd1393964494, `RNS_PRIME_BITS'd1467479091, `RNS_PRIME_BITS'd93058891, `RNS_PRIME_BITS'd377262823, `RNS_PRIME_BITS'd796221513, `RNS_PRIME_BITS'd587837481, `RNS_PRIME_BITS'd268706943},
    '{`RNS_PRIME_BITS'd2113944841, `RNS_PRIME_BITS'd1971650828, `RNS_PRIME_BITS'd624065401, `RNS_PRIME_BITS'd271566352, `RNS_PRIME_BITS'd1051786406, `RNS_PRIME_BITS'd1848214536, `RNS_PRIME_BITS'd531632460, `RNS_PRIME_BITS'd1716054783, `RNS_PRIME_BITS'd1013332612, `RNS_PRIME_BITS'd8508976, `RNS_PRIME_BITS'd1812041745, `RNS_PRIME_BITS'd1294117088, `RNS_PRIME_BITS'd602291994, `RNS_PRIME_BITS'd1262688818, `RNS_PRIME_BITS'd1869509655, `RNS_PRIME_BITS'd1960509946, `RNS_PRIME_BITS'd1714061643, `RNS_PRIME_BITS'd2035490122, `RNS_PRIME_BITS'd1805451593, `RNS_PRIME_BITS'd480486321, `RNS_PRIME_BITS'd1348869430, `RNS_PRIME_BITS'd210379497, `RNS_PRIME_BITS'd219162379, `RNS_PRIME_BITS'd1148913620, `RNS_PRIME_BITS'd305150941, `RNS_PRIME_BITS'd1397283234, `RNS_PRIME_BITS'd2006122730, `RNS_PRIME_BITS'd171919279, `RNS_PRIME_BITS'd536327602, `RNS_PRIME_BITS'd1329388365, `RNS_PRIME_BITS'd1974613206, `RNS_PRIME_BITS'd676472523, `RNS_PRIME_BITS'd516841753, `RNS_PRIME_BITS'd1635059530, `RNS_PRIME_BITS'd206088228, `RNS_PRIME_BITS'd1978964303, `RNS_PRIME_BITS'd530277962, `RNS_PRIME_BITS'd518870814, `RNS_PRIME_BITS'd1100050078, `RNS_PRIME_BITS'd1223389601, `RNS_PRIME_BITS'd232806416, `RNS_PRIME_BITS'd2109715245, `RNS_PRIME_BITS'd1009260182, `RNS_PRIME_BITS'd1880309153, `RNS_PRIME_BITS'd255993234, `RNS_PRIME_BITS'd73643954, `RNS_PRIME_BITS'd365178688, `RNS_PRIME_BITS'd1687722945, `RNS_PRIME_BITS'd1194694038, `RNS_PRIME_BITS'd1089849203, `RNS_PRIME_BITS'd710114276, `RNS_PRIME_BITS'd586395470, `RNS_PRIME_BITS'd533019697, `RNS_PRIME_BITS'd785507157, `RNS_PRIME_BITS'd944229547, `RNS_PRIME_BITS'd621626299, `RNS_PRIME_BITS'd282182630, `RNS_PRIME_BITS'd1181715581, `RNS_PRIME_BITS'd233193577, `RNS_PRIME_BITS'd1167177632, `RNS_PRIME_BITS'd327707007, `RNS_PRIME_BITS'd1982229971, `RNS_PRIME_BITS'd614945244, `RNS_PRIME_BITS'd1143589008},
    '{`RNS_PRIME_BITS'd2113947613, `RNS_PRIME_BITS'd681353102, `RNS_PRIME_BITS'd1214822842, `RNS_PRIME_BITS'd661265117, `RNS_PRIME_BITS'd595850019, `RNS_PRIME_BITS'd647462316, `RNS_PRIME_BITS'd621807479, `RNS_PRIME_BITS'd2086146408, `RNS_PRIME_BITS'd21134795, `RNS_PRIME_BITS'd1095737960, `RNS_PRIME_BITS'd1659943279, `RNS_PRIME_BITS'd818892796, `RNS_PRIME_BITS'd1131234638, `RNS_PRIME_BITS'd737003659, `RNS_PRIME_BITS'd152293315, `RNS_PRIME_BITS'd712173292, `RNS_PRIME_BITS'd840211036, `RNS_PRIME_BITS'd701151613, `RNS_PRIME_BITS'd1118340653, `RNS_PRIME_BITS'd2008388677, `RNS_PRIME_BITS'd901615418, `RNS_PRIME_BITS'd1631682801, `RNS_PRIME_BITS'd894989546, `RNS_PRIME_BITS'd1219619620, `RNS_PRIME_BITS'd181570311, `RNS_PRIME_BITS'd865222540, `RNS_PRIME_BITS'd1450038462, `RNS_PRIME_BITS'd1234398263, `RNS_PRIME_BITS'd823293093, `RNS_PRIME_BITS'd1985363596, `RNS_PRIME_BITS'd818331108, `RNS_PRIME_BITS'd1561855482, `RNS_PRIME_BITS'd1162473475, `RNS_PRIME_BITS'd679665385, `RNS_PRIME_BITS'd151684780, `RNS_PRIME_BITS'd189652214, `RNS_PRIME_BITS'd368403599, `RNS_PRIME_BITS'd1529671476, `RNS_PRIME_BITS'd1835710782, `RNS_PRIME_BITS'd809821929, `RNS_PRIME_BITS'd1467187245, `RNS_PRIME_BITS'd534996762, `RNS_PRIME_BITS'd562322150, `RNS_PRIME_BITS'd2032895388, `RNS_PRIME_BITS'd791949256, `RNS_PRIME_BITS'd1077481907, `RNS_PRIME_BITS'd1194674271, `RNS_PRIME_BITS'd381452777, `RNS_PRIME_BITS'd2104040240, `RNS_PRIME_BITS'd197504372, `RNS_PRIME_BITS'd945201478, `RNS_PRIME_BITS'd1372404310, `RNS_PRIME_BITS'd1194991604, `RNS_PRIME_BITS'd1695765452, `RNS_PRIME_BITS'd1967628692, `RNS_PRIME_BITS'd113472302, `RNS_PRIME_BITS'd367143186, `RNS_PRIME_BITS'd113949623, `RNS_PRIME_BITS'd1307104724, `RNS_PRIME_BITS'd1811708202, `RNS_PRIME_BITS'd936229520, `RNS_PRIME_BITS'd118485329, `RNS_PRIME_BITS'd733045511, `RNS_PRIME_BITS'd91268120}
};

parameter Ba_BASIS_poly twist_factor_ba   = '{
    '{`RNS_PRIME_BITS'd1, `RNS_PRIME_BITS'd408088301, `RNS_PRIME_BITS'd545722081, `RNS_PRIME_BITS'd2013316613, `RNS_PRIME_BITS'd1321642193, `RNS_PRIME_BITS'd321959319, `RNS_PRIME_BITS'd1021511790, `RNS_PRIME_BITS'd895733675, `RNS_PRIME_BITS'd1907272939, `RNS_PRIME_BITS'd1047887518, `RNS_PRIME_BITS'd130472541, `RNS_PRIME_BITS'd849014309, `RNS_PRIME_BITS'd1383024311, `RNS_PRIME_BITS'd2051297149, `RNS_PRIME_BITS'd572408039, `RNS_PRIME_BITS'd708487692, `RNS_PRIME_BITS'd1187016878, `RNS_PRIME_BITS'd1217688897, `RNS_PRIME_BITS'd1748729974, `RNS_PRIME_BITS'd1671387385, `RNS_PRIME_BITS'd2040483268, `RNS_PRIME_BITS'd985132875, `RNS_PRIME_BITS'd1013309155, `RNS_PRIME_BITS'd1103304400, `RNS_PRIME_BITS'd70525087, `RNS_PRIME_BITS'd1280246740, `RNS_PRIME_BITS'd1423738182, `RNS_PRIME_BITS'd2108544873, `RNS_PRIME_BITS'd1332271570, `RNS_PRIME_BITS'd1752678097, `RNS_PRIME_BITS'd658442757, `RNS_PRIME_BITS'd427090976, `RNS_PRIME_BITS'd1656931938, `RNS_PRIME_BITS'd828187205, `RNS_PRIME_BITS'd863028180, `RNS_PRIME_BITS'd1908486966, `RNS_PRIME_BITS'd61269856, `RNS_PRIME_BITS'd1612421805, `RNS_PRIME_BITS'd1825676708, `RNS_PRIME_BITS'd1310355683, `RNS_PRIME_BITS'd99928383, `RNS_PRIME_BITS'd1003955160, `RNS_PRIME_BITS'd1348001053, `RNS_PRIME_BITS'd819422651, `RNS_PRIME_BITS'd1070648195, `RNS_PRIME_BITS'd1226417430, `RNS_PRIME_BITS'd1453801843, `RNS_PRIME_BITS'd997812037, `RNS_PRIME_BITS'd163057938, `RNS_PRIME_BITS'd583652742, `RNS_PRIME_BITS'd1898138826, `RNS_PRIME_BITS'd1278600277, `RNS_PRIME_BITS'd1437033183, `RNS_PRIME_BITS'd2058685992, `RNS_PRIME_BITS'd2047246327, `RNS_PRIME_BITS'd2003019592, `RNS_PRIME_BITS'd608435798, `RNS_PRIME_BITS'd843307226, `RNS_PRIME_BITS'd881750696, `RNS_PRIME_BITS'd52620857, `RNS_PRIME_BITS'd1434548924, `RNS_PRIME_BITS'd618722642, `RNS_PRIME_BITS'd1713622070, `RNS_PRIME_BITS'd2138310495}
};

parameter Ba_BASIS_poly untwist_factor_ba = '{
    '{`RNS_PRIME_BITS'd2113948747, `RNS_PRIME_BITS'd1006785901, `RNS_PRIME_BITS'd1785180724, `RNS_PRIME_BITS'd594317815, `RNS_PRIME_BITS'd1990869694, `RNS_PRIME_BITS'd1911798094, `RNS_PRIME_BITS'd1328412326, `RNS_PRIME_BITS'd859246617, `RNS_PRIME_BITS'd728697515, `RNS_PRIME_BITS'd237140755, `RNS_PRIME_BITS'd1813522587, `RNS_PRIME_BITS'd1310022712, `RNS_PRIME_BITS'd1017743359, `RNS_PRIME_BITS'd684671453, `RNS_PRIME_BITS'd305889001, `RNS_PRIME_BITS'd192208878, `RNS_PRIME_BITS'd601437576, `RNS_PRIME_BITS'd152182897, `RNS_PRIME_BITS'd1688576189, `RNS_PRIME_BITS'd719041552, `RNS_PRIME_BITS'd83935348, `RNS_PRIME_BITS'd1966926300, `RNS_PRIME_BITS'd952025002, `RNS_PRIME_BITS'd789627009, `RNS_PRIME_BITS'd2112387366, `RNS_PRIME_BITS'd1153941663, `RNS_PRIME_BITS'd1179444514, `RNS_PRIME_BITS'd1484769300, `RNS_PRIME_BITS'd1072794403, `RNS_PRIME_BITS'd1782135960, `RNS_PRIME_BITS'd657610025, `RNS_PRIME_BITS'd154833285, `RNS_PRIME_BITS'd1114971667, `RNS_PRIME_BITS'd1067078448, `RNS_PRIME_BITS'd157485542, `RNS_PRIME_BITS'd543045019, `RNS_PRIME_BITS'd583168613, `RNS_PRIME_BITS'd1342798409, `RNS_PRIME_BITS'd179082543, `RNS_PRIME_BITS'd651090985, `RNS_PRIME_BITS'd1039095048, `RNS_PRIME_BITS'd519636741, `RNS_PRIME_BITS'd1158583015, `RNS_PRIME_BITS'd353709461, `RNS_PRIME_BITS'd102336417, `RNS_PRIME_BITS'd1886504867, `RNS_PRIME_BITS'd1784632163, `RNS_PRIME_BITS'd14528353, `RNS_PRIME_BITS'd1524970994, `RNS_PRIME_BITS'd391586784, `RNS_PRIME_BITS'd1299691063, `RNS_PRIME_BITS'd2014787745, `RNS_PRIME_BITS'd1823901056, `RNS_PRIME_BITS'd1228259606, `RNS_PRIME_BITS'd971048885, `RNS_PRIME_BITS'd990269018, `RNS_PRIME_BITS'd1413052767, `RNS_PRIME_BITS'd1428858068, `RNS_PRIME_BITS'd1527557011, `RNS_PRIME_BITS'd766728452, `RNS_PRIME_BITS'd549779955, `RNS_PRIME_BITS'd136315638, `RNS_PRIME_BITS'd1098779579, `RNS_PRIME_BITS'd1503587011}
};

// fastBConv precalculated inverses
parameter rns_residue_t z_MOD_q[`q_BASIS_LEN] = '{`RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd1340848717, `RNS_PRIME_BITS'd1950706637, `RNS_PRIME_BITS'd136505383, `RNS_PRIME_BITS'd1261863396, `RNS_PRIME_BITS'd490720514, `RNS_PRIME_BITS'd2048232271, `RNS_PRIME_BITS'd561180295, `RNS_PRIME_BITS'd2064343317, `RNS_PRIME_BITS'd1284162414, `RNS_PRIME_BITS'd426116969};
parameter rns_residue_t z_MOD_B[`B_BASIS_LEN] = '{`RNS_PRIME_BITS'd400603566, `RNS_PRIME_BITS'd1317047788, `RNS_PRIME_BITS'd1877527982, `RNS_PRIME_BITS'd816591707, `RNS_PRIME_BITS'd1500256234, `RNS_PRIME_BITS'd8640588, `RNS_PRIME_BITS'd1509953789, `RNS_PRIME_BITS'd1256593971, `RNS_PRIME_BITS'd1660146682, `RNS_PRIME_BITS'd390117507};
parameter rns_residue_t y_q_TO_qBBa[`qBBa_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd122, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1514938357, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1663002026, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1202970911, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1254269319, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd15070697, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd93592423, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd345241794, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd126359634, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1571891470, `RNS_PRIME_BITS'd0 },
'{ `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd0, `RNS_PRIME_BITS'd1004678308 },
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};
parameter rns_residue_t y_B_TO_Ba[`Ba_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd33728781, `RNS_PRIME_BITS'd1756228743, `RNS_PRIME_BITS'd487215260, `RNS_PRIME_BITS'd501135696, `RNS_PRIME_BITS'd459470026, `RNS_PRIME_BITS'd1877657833, `RNS_PRIME_BITS'd50297305, `RNS_PRIME_BITS'd56214635, `RNS_PRIME_BITS'd1200871039, `RNS_PRIME_BITS'd1750218591 }
};
parameter rns_residue_t y_B_TO_q[`q_BASIS_LEN][`B_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd158, `RNS_PRIME_BITS'd24, `RNS_PRIME_BITS'd203, `RNS_PRIME_BITS'd10, `RNS_PRIME_BITS'd55, `RNS_PRIME_BITS'd218, `RNS_PRIME_BITS'd198, `RNS_PRIME_BITS'd87, `RNS_PRIME_BITS'd62, `RNS_PRIME_BITS'd92 },
'{ `RNS_PRIME_BITS'd1219156511, `RNS_PRIME_BITS'd1608499681, `RNS_PRIME_BITS'd371154937, `RNS_PRIME_BITS'd924754142, `RNS_PRIME_BITS'd2003633539, `RNS_PRIME_BITS'd627440795, `RNS_PRIME_BITS'd1066486116, `RNS_PRIME_BITS'd1296251710, `RNS_PRIME_BITS'd1679092476, `RNS_PRIME_BITS'd772683368 },
'{ `RNS_PRIME_BITS'd1367502590, `RNS_PRIME_BITS'd1413619003, `RNS_PRIME_BITS'd1604587363, `RNS_PRIME_BITS'd796115568, `RNS_PRIME_BITS'd154115966, `RNS_PRIME_BITS'd287007179, `RNS_PRIME_BITS'd457558717, `RNS_PRIME_BITS'd43558045, `RNS_PRIME_BITS'd1825868505, `RNS_PRIME_BITS'd2117666329 },
'{ `RNS_PRIME_BITS'd488607457, `RNS_PRIME_BITS'd725589953, `RNS_PRIME_BITS'd166254356, `RNS_PRIME_BITS'd1679376923, `RNS_PRIME_BITS'd375851890, `RNS_PRIME_BITS'd962572449, `RNS_PRIME_BITS'd40302594, `RNS_PRIME_BITS'd37730088, `RNS_PRIME_BITS'd1726493613, `RNS_PRIME_BITS'd1162981935 },
'{ `RNS_PRIME_BITS'd317361695, `RNS_PRIME_BITS'd1920884754, `RNS_PRIME_BITS'd1303976625, `RNS_PRIME_BITS'd107931280, `RNS_PRIME_BITS'd1804980561, `RNS_PRIME_BITS'd1467513527, `RNS_PRIME_BITS'd1597511531, `RNS_PRIME_BITS'd1771541117, `RNS_PRIME_BITS'd2104139963, `RNS_PRIME_BITS'd695454200 },
'{ `RNS_PRIME_BITS'd875545508, `RNS_PRIME_BITS'd1106807570, `RNS_PRIME_BITS'd531200008, `RNS_PRIME_BITS'd656659131, `RNS_PRIME_BITS'd318605813, `RNS_PRIME_BITS'd571007940, `RNS_PRIME_BITS'd1098654767, `RNS_PRIME_BITS'd1477330056, `RNS_PRIME_BITS'd1569331694, `RNS_PRIME_BITS'd503094350 },
'{ `RNS_PRIME_BITS'd2014745094, `RNS_PRIME_BITS'd1203280856, `RNS_PRIME_BITS'd1874657457, `RNS_PRIME_BITS'd664236066, `RNS_PRIME_BITS'd1343163396, `RNS_PRIME_BITS'd349851856, `RNS_PRIME_BITS'd327986115, `RNS_PRIME_BITS'd1527009020, `RNS_PRIME_BITS'd1664893238, `RNS_PRIME_BITS'd2028124638 },
'{ `RNS_PRIME_BITS'd17214643, `RNS_PRIME_BITS'd1528026480, `RNS_PRIME_BITS'd707649348, `RNS_PRIME_BITS'd506168135, `RNS_PRIME_BITS'd623405378, `RNS_PRIME_BITS'd1082352090, `RNS_PRIME_BITS'd1990243254, `RNS_PRIME_BITS'd747636934, `RNS_PRIME_BITS'd1326828836, `RNS_PRIME_BITS'd1378524818 },
'{ `RNS_PRIME_BITS'd1873007184, `RNS_PRIME_BITS'd1982800586, `RNS_PRIME_BITS'd1616965474, `RNS_PRIME_BITS'd936503592, `RNS_PRIME_BITS'd265687623, `RNS_PRIME_BITS'd555195787, `RNS_PRIME_BITS'd703316243, `RNS_PRIME_BITS'd1230764655, `RNS_PRIME_BITS'd220437154, `RNS_PRIME_BITS'd1158294204 },
'{ `RNS_PRIME_BITS'd1171115647, `RNS_PRIME_BITS'd1636056387, `RNS_PRIME_BITS'd89367338, `RNS_PRIME_BITS'd1569217605, `RNS_PRIME_BITS'd148010597, `RNS_PRIME_BITS'd552135592, `RNS_PRIME_BITS'd1046145070, `RNS_PRIME_BITS'd1622489461, `RNS_PRIME_BITS'd627687042, `RNS_PRIME_BITS'd765167266 },
'{ `RNS_PRIME_BITS'd1810327907, `RNS_PRIME_BITS'd659636710, `RNS_PRIME_BITS'd527709368, `RNS_PRIME_BITS'd1981502868, `RNS_PRIME_BITS'd395782026, `RNS_PRIME_BITS'd1625981468, `RNS_PRIME_BITS'd263854684, `RNS_PRIME_BITS'd1651540472, `RNS_PRIME_BITS'd1368489211, `RNS_PRIME_BITS'd1257824607 }
};
parameter rns_residue_t y_q_TO_BBa[`B_BASIS_LEN +`Ba_BASIS_LEN][`q_BASIS_LEN] = '{
'{ `RNS_PRIME_BITS'd891343375, `RNS_PRIME_BITS'd600171900, `RNS_PRIME_BITS'd1603585445, `RNS_PRIME_BITS'd690197685, `RNS_PRIME_BITS'd1648248626, `RNS_PRIME_BITS'd920263580, `RNS_PRIME_BITS'd1150329475, `RNS_PRIME_BITS'd651747908, `RNS_PRIME_BITS'd613298131, `RNS_PRIME_BITS'd1031542234, `RNS_PRIME_BITS'd1378497069 },
'{ `RNS_PRIME_BITS'd288677486, `RNS_PRIME_BITS'd614060226, `RNS_PRIME_BITS'd1033890425, `RNS_PRIME_BITS'd815724763, `RNS_PRIME_BITS'd49469365, `RNS_PRIME_BITS'd62061567, `RNS_PRIME_BITS'd1147950992, `RNS_PRIME_BITS'd795171146, `RNS_PRIME_BITS'd995533003, `RNS_PRIME_BITS'd2003251247, `RNS_PRIME_BITS'd821322321 },
'{ `RNS_PRIME_BITS'd734467932, `RNS_PRIME_BITS'd2095955847, `RNS_PRIME_BITS'd1604696199, `RNS_PRIME_BITS'd1265905361, `RNS_PRIME_BITS'd776440121, `RNS_PRIME_BITS'd519547542, `RNS_PRIME_BITS'd45231263, `RNS_PRIME_BITS'd1685031663, `RNS_PRIME_BITS'd1689775415, `RNS_PRIME_BITS'd181826090, `RNS_PRIME_BITS'd290921744 },
'{ `RNS_PRIME_BITS'd1332295875, `RNS_PRIME_BITS'd390583230, `RNS_PRIME_BITS'd882270282, `RNS_PRIME_BITS'd1725949935, `RNS_PRIME_BITS'd1081809067, `RNS_PRIME_BITS'd546816522, `RNS_PRIME_BITS'd1653899216, `RNS_PRIME_BITS'd510872414, `RNS_PRIME_BITS'd1093633044, `RNS_PRIME_BITS'd766308621, `RNS_PRIME_BITS'd666708590 },
'{ `RNS_PRIME_BITS'd1758033742, `RNS_PRIME_BITS'd1578919505, `RNS_PRIME_BITS'd1865398228, `RNS_PRIME_BITS'd1843698483, `RNS_PRIME_BITS'd1254072644, `RNS_PRIME_BITS'd1055534362, `RNS_PRIME_BITS'd515625118, `RNS_PRIME_BITS'd1583301543, `RNS_PRIME_BITS'd62842952, `RNS_PRIME_BITS'd441768689, `RNS_PRIME_BITS'd962688836 },
'{ `RNS_PRIME_BITS'd2041418022, `RNS_PRIME_BITS'd978801754, `RNS_PRIME_BITS'd9263828, `RNS_PRIME_BITS'd9925530, `RNS_PRIME_BITS'd2028173586, `RNS_PRIME_BITS'd1319254538, `RNS_PRIME_BITS'd13895742, `RNS_PRIME_BITS'd1091117518, `RNS_PRIME_BITS'd516953991, `RNS_PRIME_BITS'd23821272, `RNS_PRIME_BITS'd1849178827 },
'{ `RNS_PRIME_BITS'd674062587, `RNS_PRIME_BITS'd1070000367, `RNS_PRIME_BITS'd487315302, `RNS_PRIME_BITS'd422927882, `RNS_PRIME_BITS'd82215022, `RNS_PRIME_BITS'd745172920, `RNS_PRIME_BITS'd1118399886, `RNS_PRIME_BITS'd715724108, `RNS_PRIME_BITS'd1065293916, `RNS_PRIME_BITS'd1670130875, `RNS_PRIME_BITS'd1097422041 },
'{ `RNS_PRIME_BITS'd1930327791, `RNS_PRIME_BITS'd564237487, `RNS_PRIME_BITS'd559689642, `RNS_PRIME_BITS'd1326477308, `RNS_PRIME_BITS'd1225283679, `RNS_PRIME_BITS'd1578340088, `RNS_PRIME_BITS'd2026697752, `RNS_PRIME_BITS'd668775664, `RNS_PRIME_BITS'd1054570822, `RNS_PRIME_BITS'd1243754760, `RNS_PRIME_BITS'd1554693450 },
'{ `RNS_PRIME_BITS'd1406620872, `RNS_PRIME_BITS'd1296310582, `RNS_PRIME_BITS'd147593610, `RNS_PRIME_BITS'd1963782344, `RNS_PRIME_BITS'd1354015071, `RNS_PRIME_BITS'd764583033, `RNS_PRIME_BITS'd196791480, `RNS_PRIME_BITS'd557451634, `RNS_PRIME_BITS'd1657227705, `RNS_PRIME_BITS'd1098441865, `RNS_PRIME_BITS'd1236628959 },
'{ `RNS_PRIME_BITS'd429127205, `RNS_PRIME_BITS'd1864444482, `RNS_PRIME_BITS'd1782848107, `RNS_PRIME_BITS'd566685585, `RNS_PRIME_BITS'd570883256, `RNS_PRIME_BITS'd2056772120, `RNS_PRIME_BITS'd2068655427, `RNS_PRIME_BITS'd1200192863, `RNS_PRIME_BITS'd894112574, `RNS_PRIME_BITS'd959905133, `RNS_PRIME_BITS'd327297224 },
'{ `RNS_PRIME_BITS'd843366860, `RNS_PRIME_BITS'd345904837, `RNS_PRIME_BITS'd1789186737, `RNS_PRIME_BITS'd1226376188, `RNS_PRIME_BITS'd1294545564, `RNS_PRIME_BITS'd1863458861, `RNS_PRIME_BITS'd49787340, `RNS_PRIME_BITS'd1749629066, `RNS_PRIME_BITS'd919244077, `RNS_PRIME_BITS'd1941818346, `RNS_PRIME_BITS'd1328125817 }
};

// mod switch from qBBa to BBa (precalculated finv constants)
parameter rns_residue_t qinv_MOD_BBa[`BBa_BASIS_LEN] = '{`RNS_PRIME_BITS'd1685594561, `RNS_PRIME_BITS'd1127635584, `RNS_PRIME_BITS'd1831397647, `RNS_PRIME_BITS'd1452117633, `RNS_PRIME_BITS'd1199363927, `RNS_PRIME_BITS'd1821452128, `RNS_PRIME_BITS'd953961963, `RNS_PRIME_BITS'd7988901, `RNS_PRIME_BITS'd645938236, `RNS_PRIME_BITS'd541478048, `RNS_PRIME_BITS'd433791376};

`define REG_NPOLY 12// how many polynomials can the register file store

// ---------------------------
// Operation/Control Types
// ---------------------------

// If you ever want to explicitly tag A vs B in code:
typedef enum logic [0:0] {
  POLY_A = 1'b0,
  POLY_B = 1'b1
} poly_sel_e;

typedef enum logic [1:0] {
    NO_OP,
    OP_CT_CT_ADD,
    OP_CT_PT_ADD,
    OP_CT_PT_MUL
} op_e;

typedef struct packed {
  op_e                          mode;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx1_b;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_a;
  logic [$clog2(`REG_NPOLY)-1:0]      idx2_b;
  logic [$clog2(`REG_NPOLY)-1:0]      out_a;
  logic [$clog2(`REG_NPOLY)-1:0]      out_b;
} operation;


`endif
