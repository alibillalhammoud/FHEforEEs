`include "types.svh"

`ifndef CTEXAMPLES_SVH
`define CTEXAMPLES_SVH


const rns_residue_t A1__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{82, 1007849158, 344623035, 974553355, 252232956, 1591552870, 1997619035, 168382023, 978517921, 225318580, 108420664},
    '{205, 1228814435, 151413131, 2050222428, 1413564231, 439481772, 444027837, 985258507, 583611165, 2035531980, 386692334},
    '{136, 128486397, 1816285854, 863587800, 267914966, 1697223387, 1705853764, 775183607, 1128390963, 380101658, 1930921843},
    '{232, 135710087, 1425278094, 1559673485, 176413468, 136727317, 1385941432, 1576270542, 71341352, 2081847665, 475256072},
    '{50, 717104875, 2051774700, 368829184, 6013804, 383335523, 965384056, 1828281782, 407992677, 839636323, 1460582641},
    '{142, 238512322, 2095782834, 1926466631, 348242689, 1452579508, 2076181866, 946667019, 248454984, 2108208234, 1417627426},
    '{253, 2072819984, 1872956090, 534439250, 461321156, 1648784831, 1125878975, 562094147, 1584847967, 2030964712, 362752790},
    '{234, 1457932833, 1554698931, 136975177, 1209489831, 1234868194, 1474258431, 1725337056, 1411870778, 2058986111, 157537645},
    '{211, 771191296, 1929166853, 220566812, 1515595715, 1047050759, 262115771, 1924947401, 512489747, 580532616, 1945613104},
    '{228, 1929758221, 1996127246, 937804862, 1288253295, 1076311145, 144918156, 1842504095, 1278919215, 556241807, 100699118},
    '{234, 1661095827, 20449632, 1121730000, 361938300, 1772251391, 254315466, 438135027, 876666992, 798295796, 1458298158},
    '{68, 916253055, 108274752, 1697816182, 903388280, 1716351348, 547309949, 1021283545, 1558943094, 38353636, 292512990},
    '{218, 1132664726, 1787992750, 1099387607, 1306070432, 1905096779, 1508222052, 325083905, 3522864, 959819657, 852525655},
    '{46, 487660555, 1061893582, 1972644058, 812108973, 1827722725, 285697904, 754991627, 69473664, 1068745859, 877540689},
    '{41, 1516766091, 1468304672, 792042504, 665252307, 1182398267, 1478596903, 1625334052, 1204101513, 1517514452, 1852392826},
    '{33, 235675091, 1215871282, 1745394775, 547832513, 832031840, 1084796080, 1494828160, 917052292, 1092506897, 1715992980},
    '{171, 1277622228, 687833643, 126756375, 765208504, 1634973533, 114865935, 491511062, 1938597003, 715389181, 1443341153},
    '{6, 1825586477, 1396430759, 1303407128, 1445475149, 424619735, 41354298, 1409837468, 278181591, 1819301706, 1848035921},
    '{50, 1904686822, 1106318626, 644769538, 923417179, 1061536840, 206347908, 960907922, 2014200918, 1799695897, 184868460},
    '{2, 1660605546, 1932790523, 107468360, 1475935526, 2137031813, 1842075581, 1534159273, 1414891420, 114674984, 422161172},
    '{117, 1467716298, 1845758024, 2027318364, 1497830248, 1322321168, 1937021108, 58754948, 2075407172, 983943721, 2147117881},
    '{245, 2014655720, 1862208197, 1311559924, 1955877019, 2076220394, 257564127, 565055248, 1143569118, 791472279, 927992919},
    '{3, 1680150016, 1828982382, 250397076, 767075907, 1216694894, 1666228359, 1911095743, 947926127, 69398065, 147306452},
    '{57, 929720665, 1370616561, 1312952281, 1642055929, 1027913888, 1836041565, 812388307, 1235506155, 1868402086, 197841319},
    '{136, 828673995, 575270028, 620510798, 308787199, 1057096300, 61639648, 1980586176, 2144543143, 1035521899, 1481261841},
    '{232, 1869944373, 1813643879, 1870421688, 1548197755, 1032972630, 1961780163, 206032257, 341345352, 1296559053, 1100192790},
    '{82, 1671046886, 779176347, 395545305, 548519104, 1521713106, 1778166872, 1992360836, 307943512, 1858486778, 1217376535},
    '{104, 77607433, 445781670, 362973800, 2135267821, 762068841, 381804377, 1356500139, 1620634429, 846861628, 106730909},
    '{177, 322709120, 834254757, 393772305, 633431033, 1242279121, 583416946, 609475388, 903262245, 756641082, 236176371},
    '{31, 448215137, 901976536, 445651178, 173840560, 378485855, 1170893215, 1404566493, 1110642524, 366040601, 357099177},
    '{137, 2067638453, 1373132689, 773754097, 1816808974, 717957840, 1775229345, 333239654, 199427305, 1605368013, 946081369},
    '{168, 762782950, 1381901223, 786873016, 451947566, 71222797, 1750410703, 561271880, 402400139, 822622409, 1215563929},
    '{48, 1894558169, 1252004129, 116503006, 752064863, 218438491, 603153407, 1408479531, 814442837, 1190173409, 2137012790},
    '{181, 1366303369, 9501924, 1040884399, 402384571, 1181165213, 1573770178, 1405940624, 1024760168, 1506088651, 1013324149},
    '{101, 1144638401, 3893692, 1435611144, 554819808, 1532223950, 594106318, 772678882, 305693585, 2109818209, 980397734},
    '{219, 710389119, 381253997, 930727903, 1386770720, 891839277, 137013315, 2077681754, 146278937, 883007174, 152000087},
    '{165, 682581400, 1455981910, 878917060, 2041288751, 255425535, 423747580, 1624241031, 163998385, 1049135090, 252484763},
    '{217, 1397784951, 1865708240, 2003438866, 1733411078, 1002091085, 1221828305, 1999633365, 876370933, 1885910635, 2095966213},
    '{4, 1384564752, 433472788, 665425110, 1773817788, 213524890, 1659723709, 1906464361, 1552802447, 2049845174, 1300791096},
    '{52, 338600753, 1538317438, 1105809867, 819333801, 441715862, 1213047921, 1804074273, 549432341, 1371046953, 1519781316},
    '{79, 2129008001, 1965939120, 1344460707, 1017466165, 540703789, 615494018, 590648200, 1184685854, 1020954333, 544490801},
    '{209, 1439719799, 557730061, 163664946, 2060177819, 1658964647, 102829226, 23132681, 842827861, 67300044, 1916779228},
    '{83, 216832388, 1499638702, 215052704, 889904893, 992089543, 1968596455, 1877331516, 1711973714, 1056600617, 1040737733},
    '{186, 1064824235, 987830523, 827448682, 1881048101, 77131150, 1431760059, 671022630, 1632059779, 147984288, 444699212},
    '{155, 446909929, 1145656905, 87751062, 651823414, 2111085037, 1283873057, 435908200, 989349162, 1066794502, 751065570},
    '{8, 2035000636, 1299571809, 397159397, 1149497610, 285868357, 860170220, 957433122, 1648166161, 1850235833, 1790613488},
    '{82, 1013199338, 1968587998, 1289695665, 296590121, 280092226, 2063421943, 901372286, 737217449, 1532531378, 1550494478},
    '{33, 299380480, 255743251, 1788013446, 2049595553, 253819890, 162154740, 928213509, 718679450, 671227245, 572242555},
    '{130, 667783287, 794056254, 39422024, 170203145, 972447735, 1332479475, 714672611, 2109603880, 571950693, 762736245},
    '{123, 1115696555, 1538380880, 1548856345, 1472321400, 1043517755, 922417491, 2049492523, 212262096, 619627638, 1503925676},
    '{28, 1777896165, 1394135005, 1526298610, 1881386209, 996757604, 1031386265, 1905368146, 130410828, 717318262, 1885797622},
    '{178, 1489514692, 399680613, 1884286346, 79271719, 1697376542, 973747397, 540796709, 2020879262, 1194089328, 673980632},
    '{182, 961661966, 1775541313, 243665668, 845308960, 1018410470, 1792340588, 2076560098, 894044508, 740049617, 442752118},
    '{119, 490495528, 218892080, 258539907, 1967225852, 657983768, 948953814, 636783003, 729293999, 814288155, 93362422},
    '{155, 1412279211, 40804773, 405570514, 1438162702, 1946144078, 330336588, 1397243825, 1449491717, 1477538017, 1177794342},
    '{138, 1110789405, 626528868, 881138703, 1933195299, 1114586919, 821409919, 130646675, 1873235257, 1690386107, 721418499},
    '{62, 1484266757, 1300731878, 1409114395, 1846628098, 980139663, 703773412, 1197908194, 626823517, 1621578307, 635217709},
    '{208, 734332099, 498345152, 692737758, 1662562743, 1541319866, 1270899383, 1458093008, 760536533, 1507237810, 1939598861},
    '{256, 2089344066, 544473085, 1714517841, 1913047875, 625018383, 1267544990, 638371721, 1705055400, 1433120257, 525740258},
    '{10, 414159494, 163452829, 2111205207, 1605954173, 976805569, 2088726651, 935565441, 80201478, 397089621, 783202583},
    '{199, 1147595380, 1641914833, 1574531044, 21766817, 1653584508, 1868863705, 1930662801, 782387793, 370535898, 1969474147},
    '{110, 338759259, 132866527, 462337302, 1810257211, 271485432, 2092074032, 1225657871, 1816845920, 241185360, 845414760},
    '{31, 1747421548, 4671678, 1007692149, 1622924542, 1657536354, 1511478571, 731731277, 767316846, 1078196739, 1471576852},
    '{16, 1786397361, 1613071122, 2113126473, 1684716348, 144713126, 1880867112, 538142292, 1997060930, 1552885288, 1889412258}
};

const rns_residue_t B1__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{164, 1112177129, 533724018, 177369642, 1679005539, 53351151, 2070494231, 1541419757, 1696370584, 347098394, 437246425},
    '{188, 1073643523, 1839593152, 1737833869, 475564003, 1170319952, 1652591677, 1893033484, 1289139608, 1822810015, 901509049},
    '{216, 1573781463, 993476669, 1507418708, 874189345, 692173683, 1932035895, 102459850, 954571405, 326083750, 1858900645},
    '{237, 642013974, 330177291, 1879332416, 427739881, 26936754, 532533065, 238101500, 353341552, 1979250593, 1650878797},
    '{202, 1535568654, 1348127997, 1184988662, 775725998, 1284421050, 1875436924, 555592031, 1809645727, 421487266, 1836811102},
    '{60, 1805432572, 1479444956, 244255772, 1224792621, 319799473, 347843552, 36778632, 675486343, 2009285989, 294120590},
    '{134, 1986164299, 1598529120, 1436650053, 1643346751, 272751406, 2007774722, 709297180, 75598111, 559874537, 2069463409},
    '{113, 1573748398, 454327867, 1498198574, 2111692289, 49349787, 1863696371, 1862307614, 695707079, 1806252203, 285885356},
    '{81, 793712966, 1379276323, 940594248, 251432029, 1054277901, 1259679507, 1875681120, 94997645, 1179282860, 1651078168},
    '{160, 1175247393, 1859984809, 1570158002, 686201950, 1310180575, 224171677, 358778910, 1044836134, 1536609293, 996445963},
    '{83, 1209786133, 120134477, 542613025, 1303774553, 1945101820, 1838674287, 2099921014, 1995139141, 216989535, 1052103704},
    '{154, 323465262, 1919920335, 2120776926, 1636300435, 1539610204, 155259356, 1954766996, 585577789, 1447080485, 623930339},
    '{114, 1317357697, 563472139, 1848835297, 1030568413, 473560243, 303622603, 258042912, 1350930065, 1206935250, 2026007439},
    '{142, 273472673, 1009731303, 1449642611, 552032416, 1095771467, 1077074838, 2009540474, 1904124801, 1728187139, 39381265},
    '{118, 114973467, 1032654111, 424623647, 622386705, 958463838, 2083997397, 463044866, 1928399823, 1147380493, 1306913884},
    '{18, 205335063, 1886108379, 417507717, 1311297209, 1761787574, 733919295, 379871043, 1672289111, 2033261301, 470497663},
    '{19, 929474100, 931895368, 1135264551, 904652826, 26041372, 1282426129, 325859245, 285135056, 1076641535, 781758219},
    '{36, 2087640943, 111135999, 603708949, 1834610488, 1555370594, 2081115710, 1997540534, 1116957688, 41882368, 829777403},
    '{200, 1137914062, 1836344919, 520131276, 38364962, 1536109202, 1684360181, 905999782, 713215539, 474109680, 37534418},
    '{64, 50724856, 441216684, 1558450073, 175251215, 1427316833, 1325475737, 1883296117, 972722946, 591159604, 1257059940},
    '{151, 1790526298, 1142469265, 846814022, 1632341827, 686687227, 1030300000, 885556595, 300196477, 2118400296, 2120870940},
    '{104, 274699927, 251379310, 1526905371, 122336813, 341917247, 1485190404, 1444780683, 1826772566, 280136859, 99978012},
    '{173, 856480771, 1599804980, 2118686351, 2092037919, 747563729, 2060261768, 1561048654, 1061630523, 1455980166, 242505756},
    '{80, 1974415339, 119315054, 1564842321, 1660438747, 1550063704, 717930394, 1211259338, 1241714250, 793254046, 846536773},
    '{228, 143359175, 172540776, 932916070, 1922634533, 1868506359, 714680181, 1074790159, 1345953700, 2128692627, 202642547},
    '{47, 1117142210, 1679150616, 528529137, 1873055888, 2015238493, 718828362, 2144090113, 676470118, 96294373, 1772680642},
    '{83, 996309165, 1207918232, 807082959, 1936000263, 751961263, 1436729800, 1193790209, 2037821185, 1037098591, 1288545473},
    '{233, 833129397, 1902828235, 930672876, 228521519, 922443346, 1348733275, 2075808, 1161009866, 1292162685, 12766119},
    '{126, 790372, 81104610, 1539322725, 707502649, 575965510, 283699902, 347711999, 1982566773, 968607687, 205361198},
    '{72, 1697214270, 2070533899, 1249720437, 1338706745, 1732282582, 250645441, 2059198498, 566771232, 1647576203, 1653833294},
    '{94, 629085881, 617284009, 1259963447, 479018809, 57176881, 406981233, 299561556, 1919910668, 837949126, 392964044},
    '{4, 1155221626, 1115962719, 1107701070, 1884712944, 1906075554, 1485486613, 11167577, 1120042162, 567908486, 224547887},
    '{82, 1965386384, 269005161, 242053564, 610786302, 1838563798, 1476567249, 2059693533, 1777827796, 670852388, 844248888},
    '{91, 1134339825, 374409068, 1712228254, 1494014663, 1111161829, 111038965, 2002186539, 1207964587, 1283198887, 307022268},
    '{6, 951055157, 1324536092, 627027283, 1306671700, 464939953, 295729341, 828055863, 1213152908, 1335574469, 1376581909},
    '{93, 1540780196, 587249532, 685733135, 1621209726, 48171582, 141561841, 1252461035, 1787854826, 960780260, 1444163481},
    '{162, 1772712583, 82039703, 348823278, 1409838555, 1534338606, 1532893202, 536058282, 1312782605, 1973604921, 702817201},
    '{127, 684799168, 810617566, 1563868314, 2132277025, 1176205618, 1291617212, 1838737579, 1344807809, 205029332, 1054039331},
    '{253, 1957191823, 713610747, 1022258107, 137282310, 1747398000, 1678452136, 1374050502, 58494819, 1920146036, 1030312991},
    '{12, 1516519767, 153726826, 481122877, 1653785398, 1746494811, 1421695236, 1121160833, 1275308650, 1539636806, 333468000},
    '{16, 10127594, 1000689174, 313552564, 676065905, 622357239, 949605324, 384385279, 39249879, 1197981334, 949137540},
    '{100, 337931369, 1883587918, 2144223165, 855614651, 1520467346, 94829642, 1404149425, 1447443133, 1153651154, 1330699206},
    '{48, 2059688593, 1667457801, 1704998216, 212898688, 1283772960, 1816058199, 1838322636, 1715861534, 1275659244, 420883517},
    '{25, 100752787, 1003691475, 1891578874, 17834090, 760348900, 1518570040, 803557864, 289166598, 1465043885, 803412714},
    '{249, 1717345784, 1366360348, 23323035, 1158294019, 1463842811, 618382164, 2089062547, 323297971, 1548543634, 984931701},
    '{63, 937164559, 2051324299, 1359881548, 1048106072, 197283873, 1088081970, 600312125, 860429775, 1631863013, 873653663},
    '{85, 199733385, 1229119, 581351261, 400306788, 1275471543, 1314617845, 871309140, 507070491, 72930676, 264662275},
    '{110, 1535323094, 2110171527, 181617893, 1240107990, 1760785827, 625690953, 918847505, 1121377264, 913794679, 176667167},
    '{228, 1524898392, 328776342, 1478926205, 638627153, 1525155906, 190214825, 939014537, 1370006499, 1472770738, 1901673828},
    '{225, 1977356419, 1416042110, 1268940098, 1599005508, 1360518251, 1852933215, 1845618624, 1221987484, 1025654898, 2022986732},
    '{16, 1924168719, 1117521149, 1349322214, 1825385249, 722760803, 1514640851, 713033627, 1186258764, 2082051839, 665342042},
    '{70, 1624957882, 1323885445, 105666162, 1300983833, 1840544033, 1383379926, 922984325, 19271487, 270741065, 432310072},
    '{153, 1783258660, 1233720022, 2057058461, 932263646, 1711607144, 922882246, 2003002430, 1659266438, 1540243119, 1212675658},
    '{10, 767797460, 449130898, 487780479, 912922911, 805659668, 1076739181, 1976663147, 102864022, 1144022461, 570311395},
    '{32, 1787518897, 2129617489, 1795316463, 1508132779, 910772726, 823915451, 1567449857, 1749834906, 1936884195, 416712942},
    '{40, 1880538070, 1797055427, 1032899401, 28386578, 933519243, 2015643943, 587367817, 575599096, 963794549, 322785847},
    '{120, 1767143481, 1171034278, 801826112, 129903151, 1285551010, 98640459, 1499448647, 213863181, 990285516, 564816723},
    '{146, 349263378, 1725167867, 294977853, 1364875384, 1630016139, 20313273, 959416456, 1023240651, 844469708, 756943719},
    '{216, 287220864, 1433201783, 1598528648, 1239915840, 940797769, 922005843, 552867908, 180967113, 1437316834, 452718313},
    '{245, 1580529675, 230279239, 743086191, 532454816, 1607468248, 966242335, 501280583, 726033383, 915813203, 1232024914},
    '{224, 755984682, 825850527, 867645482, 741438072, 1015419087, 1868974263, 1280052164, 576935286, 1803245003, 862452203},
    '{209, 195958570, 1678176313, 1768673732, 377441428, 283910164, 714687245, 1414491619, 1114772996, 2038631762, 1235495759},
    '{137, 711514740, 1837214213, 1945467505, 605421544, 558182535, 716094237, 1114379824, 271557769, 2097514290, 1782698781},
    '{200, 707719628, 988967764, 2055368146, 1745192673, 177037800, 1835330505, 1017619763, 182878640, 546019738, 357572893}
};

const rns_residue_t A2__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{36, 1340328697, 1028411192, 833505390, 508914425, 695101177, 121929651, 468190141, 158621671, 1229496176, 1922507611},
    '{227, 1897012015, 424664047, 148390489, 1660881012, 1839841661, 600890401, 111859334, 63012075, 1837715341, 2102711601},
    '{177, 952024879, 1847294303, 1024507888, 1731714129, 456798983, 398357807, 819150038, 1074871179, 1881538838, 984786775},
    '{5, 214890831, 1793609357, 293158148, 941952042, 1703338787, 477362987, 755957961, 1779634707, 886758664, 322190161},
    '{21, 2013309932, 1196272423, 1913281042, 1933756359, 1005191015, 2100169185, 186901693, 1462544178, 642790623, 150495599},
    '{101, 712620492, 253161811, 171550392, 2035805351, 2095024128, 1227883816, 575815669, 2002458832, 1563852721, 508758874},
    '{13, 832585577, 357443542, 283467771, 856202594, 1002737735, 782790808, 1985333376, 245128879, 351791664, 1185501061},
    '{7, 293386272, 1188507358, 22433621, 582320240, 2094628288, 828243241, 1318815447, 1561322294, 251856247, 586126026},
    '{111, 707227732, 2074311491, 2131174023, 567084629, 1168712801, 1143862775, 399711304, 1164710298, 237095739, 1223221511},
    '{104, 713648247, 479395508, 289517191, 270218379, 2100172118, 1611389917, 1301115129, 728629924, 1579218442, 271989711},
    '{246, 237400224, 1139042970, 282688036, 869650008, 491537767, 1441081581, 655100268, 1557975835, 1026539034, 499527145},
    '{177, 557753617, 878833429, 1373561798, 1844073307, 94445269, 2014326158, 343865196, 775191453, 1608547572, 126311803},
    '{82, 252932985, 1123198115, 896914588, 969680251, 1168800444, 1914069947, 263023560, 799316948, 352769466, 313895061},
    '{90, 1771618026, 1407987179, 1723691945, 721970711, 1012620522, 404576311, 57230767, 1868541068, 1152816320, 621194939},
    '{181, 1242370691, 1436402501, 1305837762, 1420137746, 57070319, 1789467850, 586454966, 549398473, 595211950, 74535715},
    '{59, 363925171, 1086348616, 353727616, 373279121, 518645799, 1473668681, 744013713, 629613559, 1943859100, 789731493},
    '{230, 1218992033, 2056101164, 483236890, 347881410, 718379194, 89425199, 1226296273, 721891169, 2066476512, 1804991562},
    '{136, 455237887, 1892988214, 1279868935, 603784556, 212834038, 492818166, 349005833, 856605567, 566636026, 200972298},
    '{215, 352156915, 416537380, 2057979471, 521394630, 520005871, 1371324822, 95777377, 138940384, 1847750006, 626091291},
    '{70, 1765902167, 237580393, 1583354238, 881356348, 55580668, 447871555, 495777285, 1402912932, 1589862690, 1961501413},
    '{174, 452946413, 1648354070, 1953678431, 1895756983, 327607571, 306136394, 893032770, 1339902012, 907888793, 2096271269},
    '{17, 530928021, 1045149885, 620184326, 1854123236, 164062551, 1709464154, 168182394, 334728737, 213279582, 1255432417},
    '{191, 1202546534, 1254129065, 1579796147, 1787262223, 1705922028, 508253148, 1313033174, 807185662, 259916130, 456307767},
    '{82, 34800640, 1761558539, 228331537, 1422312480, 432608989, 1148635437, 1685559959, 1710561155, 670637027, 101903952},
    '{38, 1563853717, 571201328, 245251714, 1663970889, 1902173506, 189846866, 1451639541, 1558590312, 2006475795, 731899446},
    '{181, 953006543, 1333419366, 803996697, 699638571, 1570575928, 1754980088, 706796035, 1027625782, 2133888631, 1162595841},
    '{77, 1637537897, 20482474, 889619225, 1780328347, 1517088642, 1435596795, 1930430867, 1520097171, 1029411705, 506584303},
    '{58, 1518024326, 1927616150, 1161933470, 1072463355, 2079805121, 1570064471, 149929679, 306716022, 1496495185, 1041866057},
    '{178, 1400343730, 32890735, 1645109039, 332720266, 522951379, 1266211659, 1374693309, 874681560, 204708434, 609873395},
    '{205, 2117964355, 1542791771, 259735212, 1640745609, 1283940151, 929408010, 1005391845, 295962104, 18063076, 2128075980},
    '{229, 1385643703, 726954292, 1736206351, 680972654, 1491864843, 930967383, 1412993692, 1701231324, 983954389, 775122167},
    '{242, 682683785, 1458002286, 130064439, 515229608, 240014085, 732547739, 700413047, 1405345957, 290637115, 990713641},
    '{96, 364431565, 1277017596, 1522582382, 1786416419, 861608707, 1284337464, 1071267324, 1115579539, 1943030248, 1035515045},
    '{45, 1564900277, 672953399, 533116035, 1971824569, 256140759, 550284574, 1868169509, 1949422640, 787871302, 1915179667},
    '{37, 888635231, 591286787, 2142481268, 2049260352, 1140808319, 321165315, 965976563, 1671350840, 1644418855, 1677324236},
    '{27, 1637530535, 2087681052, 1478245845, 995137290, 584188626, 1885333088, 1845090887, 428160732, 1073719221, 1448512584},
    '{253, 1749950010, 580420431, 892596393, 1019570997, 885458894, 514520152, 336938809, 1211993469, 630510729, 1561927548},
    '{236, 387697373, 1513009803, 1122647403, 423356178, 732466220, 1449223682, 855139304, 1746389734, 1042485439, 965972923},
    '{171, 1103034900, 187595593, 708552635, 195619786, 1776899433, 1897397501, 1883876023, 909312593, 1828144020, 1271430307},
    '{251, 972408796, 1667335346, 1348489626, 1422461612, 1880010760, 423612396, 507740764, 144120395, 1318962956, 619499839},
    '{16, 948585442, 13763333, 685888583, 169247853, 239620760, 725391476, 276938486, 488687644, 139413933, 556100233},
    '{112, 455635859, 2046527541, 688338515, 789628807, 776121815, 2015930360, 1039112052, 1257796053, 1363141974, 1849975529},
    '{234, 1451617879, 911347881, 830018904, 1194628656, 1301376534, 2101833799, 1029298036, 934458470, 1434806506, 50832969},
    '{132, 1923221321, 574863860, 1825964470, 1080821454, 1628149686, 1111625142, 1967290119, 963652876, 693488822, 936107445},
    '{80, 1239035345, 1396123321, 649161926, 597549788, 807581434, 1657302521, 350202451, 1469810176, 1731537838, 1473677131},
    '{225, 1927225614, 169557685, 1124531029, 645893142, 11808009, 1318488075, 399784272, 935117004, 787168005, 1311169409},
    '{179, 854068432, 320347225, 1658503202, 127165862, 578927198, 766179215, 1048877454, 941095724, 956202953, 1293147664},
    '{236, 678560121, 2109389178, 1643846849, 1393021507, 1923080752, 576549368, 1256355067, 950129201, 1498451417, 1529713522},
    '{233, 485324390, 867109936, 614876355, 813104772, 2014655754, 579028278, 637212477, 1457836900, 936084674, 1257556765},
    '{83, 1270140768, 289457166, 636248138, 420615460, 1080981210, 1715305531, 865940732, 1181573363, 85644503, 1563555965},
    '{207, 605171683, 935946349, 934562408, 692311391, 2129468798, 492377783, 370107380, 1734485218, 1953235194, 12929148},
    '{5, 845066254, 383929236, 1727537090, 524673580, 1110222294, 942316711, 710838697, 881641935, 1476192243, 1301340958},
    '{68, 523124056, 1725990315, 1802356227, 929179022, 2038391289, 763417140, 1867905882, 240396442, 1514687753, 662086514},
    '{62, 1008923926, 1712267184, 66715980, 2116786604, 1705268748, 167592567, 941595340, 2112950272, 966183466, 68405799},
    '{13, 303034312, 125642853, 1409626079, 1641311794, 943835740, 1569241352, 742445703, 1396267602, 62563416, 359370362},
    '{33, 1751464864, 523326004, 1335530113, 765454914, 1668622198, 117421188, 1924208047, 1595402938, 1870251196, 1067446201},
    '{155, 1580803029, 176956725, 1091609407, 1945581937, 1758300001, 350292717, 1114617248, 590064287, 986480542, 424378780},
    '{78, 97191010, 1363669740, 668503916, 500864865, 631297502, 1109658718, 532533810, 936353871, 936998295, 2130785219},
    '{151, 816211149, 1584074260, 1752514649, 1081668837, 474083483, 1356426305, 1086476956, 1019470604, 1037006672, 861969653},
    '{207, 1595186567, 1432874892, 1786110961, 1106254626, 1259076666, 1345402623, 119932553, 1067721364, 1368327433, 2145273054},
    '{245, 1881822655, 1087427362, 1453347102, 1629269185, 1625128790, 1399142330, 124806697, 2128518943, 835731850, 1040493708},
    '{194, 404944566, 329289509, 1147166527, 1500208368, 1075924044, 818763913, 2041605630, 33458838, 1105837464, 1741403262},
    '{149, 466007139, 2085642063, 902279933, 930674557, 843689752, 723893333, 293672503, 1732507925, 1973944467, 298255786},
    '{222, 1459654781, 914457688, 1441067476, 623050342, 1556747181, 1135592291, 1024092932, 998978140, 652166025, 1674169521}
};

const rns_residue_t B2__INPUT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{141, 819594541, 634162875, 416060616, 1154266234, 264646753, 1294044377, 950158574, 1513440422, 510797271, 489440472},
    '{207, 2099677320, 1394874675, 246679523, 147367499, 1043590720, 1582511291, 1209090269, 612566604, 738619560, 1179291959},
    '{61, 258927413, 1564853584, 2019452835, 891764881, 1359612792, 1482587554, 797572147, 477094657, 326608940, 640982479},
    '{35, 739401343, 1929523711, 1400841293, 770807617, 462147960, 1562561271, 1205264550, 1044595842, 1251653041, 552842896},
    '{88, 1247659774, 391309228, 1024538162, 1791655406, 2080402555, 1666855140, 1927242802, 1064001599, 1912116412, 1169633428},
    '{171, 1911121266, 705622760, 739670038, 909302998, 148429629, 826775930, 799157589, 878768207, 1549848747, 1203674671},
    '{39, 2063930116, 1239914681, 1512585477, 767597840, 14632487, 944296055, 794245830, 1818032962, 865915819, 1353149694},
    '{111, 2137032593, 160694811, 2042135463, 96815553, 1708371853, 2064372185, 231545039, 802166271, 1163026014, 1492809667},
    '{242, 585108949, 1637316131, 1939982992, 551816933, 601710522, 500571175, 1262582880, 2128675053, 1432919088, 71493683},
    '{88, 915546312, 1769984116, 1634450517, 1592951776, 1705215505, 1810505395, 344265869, 362893885, 773437358, 1541030359},
    '{177, 320023024, 1633694796, 1277232448, 1214945911, 1290607432, 369284065, 1622292502, 590955315, 342395329, 685387561},
    '{99, 63805056, 162020278, 1079972613, 1074912741, 320186891, 1081964390, 306135782, 748725397, 1357489484, 27601783},
    '{53, 915789616, 492156745, 1890560515, 1499642239, 738472914, 1217845942, 9513633, 302480995, 429401347, 791717471},
    '{196, 900496020, 1821279819, 370179858, 2091846939, 1733497096, 1454806985, 1911927546, 123883023, 403362424, 516266982},
    '{19, 187169408, 527880281, 1404867017, 2094678075, 235416160, 1268826050, 750702119, 1107019521, 1188608593, 1424694820},
    '{88, 1962284189, 405995601, 1860144133, 798327847, 1226026097, 183579251, 371890941, 1273651218, 1507770632, 1014435354},
    '{109, 434472083, 1195837800, 2103407449, 1965061855, 206649400, 847617629, 542249444, 398466813, 452142554, 1994865915},
    '{125, 1708886125, 21734104, 1644786707, 1133762070, 101403868, 626538050, 63595077, 401308502, 708118130, 1141714986},
    '{148, 1406336163, 917044915, 1784945458, 1807509622, 1618340064, 2056570318, 1257821790, 125273275, 940657878, 370317992},
    '{128, 2114345677, 755890230, 1785417239, 433814654, 1826163059, 1211851383, 432931089, 2102654618, 1337902534, 1923230211},
    '{238, 1764916304, 204792834, 1529220789, 754892120, 1233638851, 539059469, 950427990, 1300131394, 1911425273, 1046872352},
    '{191, 795705422, 307112129, 578197630, 790226394, 686008000, 310783029, 2105070156, 61914444, 1530203265, 343976073},
    '{130, 649620689, 290477270, 814298233, 797115476, 1141346909, 585449068, 1627518940, 207871773, 157538683, 589066518},
    '{80, 10593591, 1315039663, 1711382794, 1379485415, 1640851746, 1136932273, 423568379, 773279288, 1580401593, 990756297},
    '{123, 1037357647, 1880641985, 1815670141, 811775812, 383333173, 1925215314, 515541833, 911697722, 1950762573, 2106453894},
    '{103, 505170993, 1989781485, 1856998026, 322222697, 1120433739, 906370740, 40538344, 1546724913, 440647083, 608733416},
    '{153, 45183827, 1871540698, 2016433637, 1839729940, 1995915962, 359544319, 958241987, 1899818794, 1389431075, 514254217},
    '{102, 808516534, 288108505, 1779630902, 251205849, 1332817229, 871687549, 537877349, 1815713409, 1927809613, 2002278688},
    '{66, 1683576530, 691310118, 9759421, 315304674, 1501326164, 1343653819, 62806841, 1479987306, 408322850, 15854668},
    '{159, 685522803, 1850961960, 1338318109, 1173062036, 926763889, 219410212, 487931553, 682918181, 230619588, 1000310099},
    '{114, 1167225490, 525385688, 1745161141, 2092847354, 892798744, 1401580004, 1011219402, 465573817, 129325776, 1071014226},
    '{86, 507364865, 1563159291, 1365781818, 63469546, 1075610932, 1984736417, 1421309241, 908302736, 1952866778, 1659354016},
    '{139, 1850216090, 1876205825, 1909699202, 232283774, 315223927, 1778499475, 865164276, 1679998137, 759745973, 656494698},
    '{185, 1865733028, 667006868, 835234464, 2082753758, 760281411, 135500266, 1608769802, 514408627, 659313086, 1310779780},
    '{62, 1259530563, 476318156, 680762550, 159981766, 2033001506, 229622041, 509257478, 543362069, 103697047, 469819335},
    '{205, 1937543423, 1584544454, 1030079445, 1581533699, 287727090, 1383795100, 1357499877, 2101530144, 2109492613, 344117896},
    '{118, 1588040716, 581138958, 374659104, 1499255420, 1646577728, 1573543713, 61131976, 1228581756, 635041659, 1074368431},
    '{249, 353151116, 1901108365, 242482366, 519832031, 1392418782, 62306133, 1941131409, 1942740236, 563391762, 413079715},
    '{113, 1512092100, 1004993655, 370115863, 1875428201, 1497052943, 1585766739, 1412955168, 501302281, 702748572, 1225237193},
    '{185, 520149647, 515840591, 1498299651, 951545154, 639081141, 1059491839, 747090048, 1961143623, 400265686, 1198064782},
    '{20, 1633012320, 1899398377, 128854809, 837024261, 2036820037, 1415002192, 553634430, 2076305604, 76323298, 414637080},
    '{128, 1349680490, 1885788375, 2095417360, 1119908856, 1421065110, 1223027882, 151382369, 436880576, 1046791115, 1925704257},
    '{252, 1485058326, 163218604, 362222291, 2089249362, 1783759357, 467135732, 1902375748, 543808913, 248239272, 1626540682},
    '{37, 2071347513, 1236608507, 1737180625, 1222965153, 1691308329, 1113227519, 2001857042, 1918939872, 860140297, 1495208453},
    '{59, 1791435174, 1084854030, 621860874, 1847956270, 1433278422, 2015090342, 1140134113, 387546390, 1875855755, 1826620531},
    '{172, 1969319885, 1216157117, 730992467, 1878086538, 1020341647, 499438714, 1809855918, 1385221753, 1961683318, 37117288},
    '{56, 1239046014, 721545418, 884781362, 2141877787, 506316102, 470970923, 1225090920, 718658589, 1568470193, 1664245286},
    '{238, 2073859148, 489244135, 559889518, 1182433980, 2031475891, 42550269, 1842190454, 807987318, 269870557, 271371963},
    '{38, 984322734, 824282316, 112237508, 281203694, 1042679965, 534649879, 973730440, 587091442, 519490093, 35005606},
    '{49, 1630999126, 340531089, 1688081553, 385333044, 1878325669, 1633392792, 1807393328, 595045519, 1613425123, 219343411},
    '{23, 36729657, 1508989410, 1830400439, 82583994, 1805805965, 196658475, 278215989, 2138056788, 1724214718, 1600476637},
    '{55, 918617108, 557513931, 937998306, 157008105, 1422187120, 1083468845, 1192876938, 1579861557, 311266367, 1598272207},
    '{71, 1619949148, 1869077212, 1052858990, 1983164030, 460623130, 908142441, 435004017, 789128822, 623154567, 475302146},
    '{113, 1254656806, 939423615, 217426265, 793662265, 1438970055, 1813246673, 1760659138, 1610565970, 669839357, 515008055},
    '{207, 801292751, 125414128, 1835109919, 1590975911, 1400398193, 1787450193, 1560206241, 1107439063, 939528944, 1968363546},
    '{57, 1259738979, 661307225, 1471575602, 1224673920, 782037770, 1168354673, 1705579204, 2041561654, 412736450, 1797787300},
    '{250, 529873324, 1643627776, 176640800, 800805370, 2079567618, 1634430711, 381351272, 84392422, 1907477978, 173024401},
    '{155, 1798433420, 426691550, 2046591696, 1896915698, 1668408377, 1455614987, 122326003, 298471715, 988993182, 973820226},
    '{188, 1746944146, 689413925, 568471329, 236800199, 122139162, 1844962836, 2046340204, 1752607832, 38992540, 666891989},
    '{199, 780035199, 696210964, 2088411845, 1803926387, 1141553324, 857805867, 460171281, 1285011957, 398309669, 1149897308},
    '{131, 187755374, 290063259, 144189588, 264727077, 1186399850, 1391700886, 475214180, 103801547, 831416657, 694183002},
    '{202, 1504604023, 2051724076, 460984519, 505776639, 1257572390, 619517656, 1520366583, 588667642, 613176603, 1678891937},
    '{160, 87626930, 1428342435, 334829787, 575426957, 1135762866, 2028759844, 1925903783, 1137575117, 2035276103, 752620199},
    '{9, 1472894112, 666024268, 161246846, 770546544, 264543335, 1156921901, 347183034, 1952749082, 135120201, 816699828}
};

const rns_residue_t PLAIN__TEXT [`N_SLOTS][`q_BASIS_LEN] = '{
    '{153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153},
    '{147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147},
    '{64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64},
    '{155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155},
    '{171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171},
    '{23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23},
    '{253, 253, 253, 253, 253, 253, 253, 253, 253, 253, 253},
    '{98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98},
    '{193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193},
    '{235, 235, 235, 235, 235, 235, 235, 235, 235, 235, 235},
    '{92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92},
    '{194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194},
    '{95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95},
    '{6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6},
    '{115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115},
    '{210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210},
    '{44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44},
    '{46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46},
    '{73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73},
    '{3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3},
    '{81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81},
    '{55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55},
    '{242, 242, 242, 242, 242, 242, 242, 242, 242, 242, 242},
    '{13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13},
    '{222, 222, 222, 222, 222, 222, 222, 222, 222, 222, 222},
    '{174, 174, 174, 174, 174, 174, 174, 174, 174, 174, 174},
    '{122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122},
    '{153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153},
    '{214, 214, 214, 214, 214, 214, 214, 214, 214, 214, 214},
    '{116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116},
    '{82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82},
    '{30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30},
    '{127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127},
    '{73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73},
    '{207, 207, 207, 207, 207, 207, 207, 207, 207, 207, 207},
    '{5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5},
    '{50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50},
    '{62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62},
    '{29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29},
    '{33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33},
    '{157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157},
    '{203, 203, 203, 203, 203, 203, 203, 203, 203, 203, 203},
    '{102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102},
    '{88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88},
    '{247, 247, 247, 247, 247, 247, 247, 247, 247, 247, 247},
    '{91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91},
    '{209, 209, 209, 209, 209, 209, 209, 209, 209, 209, 209},
    '{211, 211, 211, 211, 211, 211, 211, 211, 211, 211, 211},
    '{63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63},
    '{170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170},
    '{253, 253, 253, 253, 253, 253, 253, 253, 253, 253, 253},
    '{60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60},
    '{248, 248, 248, 248, 248, 248, 248, 248, 248, 248, 248},
    '{147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147},
    '{203, 203, 203, 203, 203, 203, 203, 203, 203, 203, 203},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173},
    '{184, 184, 184, 184, 184, 184, 184, 184, 184, 184, 184},
    '{41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41},
    '{208, 208, 208, 208, 208, 208, 208, 208, 208, 208, 208},
    '{218, 218, 218, 218, 218, 218, 218, 218, 218, 218, 218},
    '{238, 238, 238, 238, 238, 238, 238, 238, 238, 238, 238},
    '{63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63},
    '{59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59}
};

const rns_residue_t PLAIN__TEXTSCALED_FORADD [`N_SLOTS][`q_BASIS_LEN] = '{
    '{162, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{236, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{173, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{228, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{116, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{99, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{235, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{162, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{151, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{238, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{74, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{96, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{189, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{171, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{199, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{233, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{180, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{187, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{89, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{190, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{252, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{233, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
};

const rns_residue_t CTCT_ADDA__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{118, 200694078, 1373034227, 1808058745, 761147381, 139167198, 2119548686, 636572164, 1137139592, 1454814756, 2030928275},
    '{175, 978342673, 576077178, 51127988, 926960186, 131836584, 1044918238, 1097117841, 646623240, 1725756120, 341911582},
    '{56, 1080511276, 1516095996, 1888095688, 1999629095, 6535521, 2104211571, 1594333645, 55771453, 114149295, 768216265},
    '{237, 350600918, 1071403290, 1852831633, 1118365510, 1840066104, 1863304419, 184738966, 1850976059, 821115128, 797446233},
    '{71, 582931030, 1100562962, 134625297, 1939770163, 1388526538, 918065240, 2015183475, 1870536855, 1482426946, 1611078240},
    '{243, 951132814, 201460484, 2098017023, 236562983, 1400116787, 1156577681, 1522482688, 103423127, 1524569754, 1926386300},
    '{9, 757921784, 82915471, 817907021, 1317523750, 504035717, 1908669783, 399937986, 1829976846, 235265175, 1548253851},
    '{241, 1751319105, 595722128, 159408798, 1791810071, 1182009633, 155013671, 896662966, 825702383, 163351157, 743663671},
    '{65, 1478419028, 1855994183, 204255906, 2082680344, 68276711, 1405978546, 177169168, 1677200045, 817628355, 1021342262},
    '{75, 495922691, 328038593, 1227322053, 1558471674, 1028996414, 1756308073, 996129687, 2007549139, 2135460249, 372688829},
    '{223, 1898496051, 1159492602, 1404418036, 1231588308, 116302309, 1695397047, 1093235295, 287152138, 1824834830, 1957825303},
    '{245, 1474006672, 987108181, 923893051, 599976530, 1810796617, 414148106, 1365148741, 186643858, 1646901208, 418824793},
    '{43, 1385597711, 763706704, 1996302195, 128265626, 926410374, 1274803998, 588107465, 802839812, 1312589123, 1166420716},
    '{136, 111794804, 322396600, 1548851074, 1534079684, 692856398, 690274215, 812222394, 1938014732, 74070978, 1498735628},
    '{222, 611653005, 757223012, 2097880266, 2085390053, 1239468586, 1120576752, 64299481, 1753499986, 2112726402, 1926928541},
    '{92, 599600262, 154735737, 2099122391, 921111634, 1350677639, 410976760, 91352336, 1546665851, 888874796, 358232120},
    '{144, 349130484, 596450646, 609993265, 1113089914, 205865878, 204291134, 1717807335, 512997483, 634374492, 1100840362},
    '{142, 133340587, 1141934812, 435791134, 2049259705, 637453773, 534172464, 1758843301, 1134787158, 238446531, 2049008219},
    '{8, 109359960, 1522856006, 555264080, 1444811809, 1581542711, 1577672730, 1056685299, 5650613, 1499954702, 810959751},
    '{72, 1279023936, 22886755, 1690822598, 209806817, 45125632, 142459135, 2029936558, 670313663, 1704537674, 236170232},
    '{34, 1920662711, 1346627933, 1833511866, 1246102174, 1649928739, 95669501, 951787718, 1267818495, 1891832514, 2095896797},
    '{5, 398099964, 759873921, 1931744250, 1662515198, 92796096, 1967028281, 733237642, 1478297855, 1004751861, 35932983},
    '{194, 735212773, 935627286, 1830193223, 406853073, 775130073, 26993506, 1076639380, 1755111789, 329314195, 603614219},
    '{139, 964521305, 984690939, 1541283818, 916883352, 1460522877, 837189001, 350458729, 798576621, 391547912, 299745271},
    '{174, 245043935, 1146471356, 865762512, 1972758088, 811782957, 251486514, 1284736180, 1555642766, 894506493, 65668934},
    '{156, 675467139, 999579084, 526933456, 100351269, 456061709, 1569272250, 912828292, 1368971134, 1282956483, 115296278},
    '{159, 1161101006, 799658821, 1285164530, 181362394, 891314899, 1066275666, 1775302166, 1828040683, 740407282, 1723960838},
    '{162, 1595631759, 225913659, 1524907270, 1060246119, 694387113, 1951868848, 1506429818, 1927350451, 195865612, 1148596966},
    '{98, 1723052850, 867145492, 2038881344, 966151299, 1765230500, 1849628605, 1984168697, 1777943805, 961349516, 846049766},
    '{236, 418695715, 297284146, 705386390, 1814586169, 1662426006, 2100301225, 262468801, 1406604628, 384103677, 337682804},
    '{109, 1305798379, 2100086981, 362475519, 350296571, 62335834, 558708727, 1746233346, 1900658629, 441831201, 1721203536},
    '{153, 1445466735, 692419348, 916937455, 967177174, 311236882, 335470441, 1261684927, 1807746096, 1113259524, 58785217},
    '{144, 111505957, 381537564, 1639085388, 390996225, 1080047198, 1887490871, 332257318, 1930022376, 985712456, 1025035482},
    '{226, 783719869, 682455323, 1574000434, 226724083, 1437305972, 2124054752, 1126620596, 826692119, 146468752, 781011463},
    '{138, 2033273632, 595180479, 1430607483, 456595103, 525545420, 915271633, 1738655445, 1977044425, 1606745863, 510229617},
    '{246, 200435877, 321450888, 261488819, 234422953, 1476027903, 2022346403, 1775283104, 574439669, 1956726395, 1600512671},
    '{161, 285047633, 2036402341, 1771513453, 913374691, 1140884429, 938267732, 1961179840, 1375991854, 1679645819, 1814412311},
    '{196, 1785482324, 1231233882, 978601340, 9282199, 1734557305, 523563986, 707283132, 475269978, 780904873, 914446783},
    '{175, 340115875, 621068381, 1373977745, 1969437574, 1990424323, 1409633209, 1642850847, 314624351, 1730497993, 424729050},
    '{46, 1311009549, 1058168623, 306814564, 94310356, 174239773, 1636660317, 164325500, 693552736, 542518708, 2139281155},
    '{95, 930109666, 1979702453, 2030349290, 1186714018, 780324549, 1340885494, 867586686, 1673373498, 1160368266, 1100591034},
    '{64, 1895355658, 456773441, 852003461, 702321569, 287599613, 2118759586, 1062244733, 2100623914, 1430442018, 1619262404},
    '{60, 1668450267, 263502422, 1045071608, 2084533549, 145979228, 1922942253, 759140015, 498941495, 343915922, 1091570702},
    '{61, 840561779, 1562694383, 505928223, 814384498, 1705280836, 395897200, 490823212, 448221966, 841473110, 1380806657},
    '{235, 1685945274, 394296065, 736912988, 1249373202, 771179622, 793687577, 786110651, 311668649, 650841139, 77250348},
    '{233, 1814742473, 1469129494, 1521690426, 1795390752, 297676366, 31170294, 1357217394, 435792476, 489912637, 954290544},
    '{4, 1867267770, 141451062, 800713938, 423755983, 859019424, 682113157, 1950249740, 1678313173, 341243130, 696149789},
    '{12, 977940601, 217648268, 1284375366, 1295132003, 29413793, 738704108, 37079039, 1668808651, 22187461, 2101956077},
    '{106, 1153107677, 1661166190, 654298379, 983307917, 839616640, 1911507753, 1351885088, 1419950091, 1508035367, 2020293010},
    '{206, 238353546, 1827838046, 37619554, 1892936860, 2124498965, 490235021, 767943718, 1393835459, 705272141, 919989288},
    '{235, 235584071, 182597193, 313376089, 426212543, 978739553, 1523764048, 127985989, 1864896046, 523062255, 1898726770},
    '{183, 187097169, 783609849, 1464338507, 603945299, 660111987, 1916064108, 1251635406, 755030508, 522790370, 1975321590},
    '{250, 1484786022, 1354047467, 2046021895, 1774487982, 909314910, 408269727, 1796976443, 1134440950, 107246169, 1104838632},
    '{181, 1499419454, 1931159264, 325255887, 1936527399, 215765667, 1116546381, 1578378343, 694753582, 1780471621, 161768221},
    '{168, 1715313523, 166447626, 1815196593, 931989439, 742492969, 1899577940, 2139689528, 698268630, 1540101433, 1537164704},
    '{171, 714770492, 1149854872, 69183887, 551165156, 635722268, 938831107, 2054854722, 1321147506, 1413146102, 1788864700},
    '{217, 917586009, 1477688603, 353238873, 1644724978, 590952815, 1054066129, 165035905, 1216887804, 460567648, 1059596489},
    '{29, 831523109, 1862014892, 1361241674, 15942551, 25130519, 233070100, 1990626818, 1696890404, 296744904, 1922891727},
    '{150, 758071438, 2128547345, 1319547561, 847231655, 1099101866, 476483294, 1724848677, 577035315, 322635728, 1387709911},
    '{217, 2009346061, 1596327721, 1749831239, 564723742, 88395386, 1286641273, 1055497994, 1147922842, 1765417054, 780983284},
    '{187, 881934258, 581858034, 880393217, 1651036002, 1131226449, 1120518034, 2055469498, 763416047, 1206267748, 862475502},
    '{47, 743703825, 462156036, 1609503829, 1162980522, 1347409476, 763349944, 1119773964, 1850304758, 1347022824, 439325669},
    '{180, 65944910, 2090313741, 1909972082, 406114042, 353739257, 87883903, 1025403780, 352334082, 904650005, 1769832638},
    '{238, 1098568365, 380044649, 1406709020, 160281633, 1701460307, 868971402, 1562235224, 848548381, 57560112, 1416089426}
};

const rns_residue_t CTCT_ADDB__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{48, 1931771670, 1167886893, 593430258, 685786716, 317997904, 1217050607, 344088794, 1062320317, 857895665, 926686897},
    '{138, 1025837066, 1086983666, 1984513392, 622931502, 66423823, 1087614967, 954634216, 1901706212, 413938374, 2080801008},
    '{20, 1832708876, 410846092, 1379386614, 1765954226, 2051786475, 1267135448, 900031997, 1431666062, 652692690, 352390771},
    '{15, 1381415317, 112216841, 1132688780, 1198547498, 489084714, 2095094336, 1443366050, 1397937394, 1083412433, 56229340},
    '{33, 635744651, 1739437225, 62041895, 419896347, 1217336756, 1394804063, 335345296, 726156637, 186112477, 858952177},
    '{231, 1569070061, 37583555, 983925810, 2134095619, 468229102, 1174619482, 835936221, 1554254550, 1411643535, 1497795261},
    '{173, 1902610638, 690959640, 801750601, 263459534, 287383893, 804582776, 1503543010, 1893631073, 1425790356, 1275120750},
    '{224, 1563297214, 615022678, 1392849108, 61022785, 1757721640, 1780580555, 2093852653, 1497873350, 821787016, 1778695023},
    '{66, 1378821915, 869108293, 733092311, 803248962, 1655988423, 1760250682, 990774463, 76182009, 464710747, 1722571851},
    '{248, 2090793705, 1482484764, 1057123590, 131668669, 867909231, 2034677072, 703044779, 1407730019, 162555450, 389983969},
    '{3, 1529809157, 1753829273, 1819845473, 371235407, 1088222403, 60470351, 1574723979, 438603767, 559384864, 1737491265},
    '{253, 387270318, 2081940613, 1053264610, 563728119, 1859797095, 1237223746, 113413241, 1334303186, 657078768, 651532122},
    '{167, 85663536, 1055628884, 1591910883, 382725595, 1212033157, 1521468545, 267556545, 1653411060, 1636336597, 670232557},
    '{81, 1173968693, 683526961, 1819822469, 496394298, 681781714, 384393822, 1773978483, 2028007824, 2131549563, 555648247},
    '{137, 302142875, 1560534392, 1829490664, 569579723, 1193879998, 1205335446, 1213746985, 887928655, 188497885, 584116351},
    '{106, 20135475, 144619819, 130166921, 2109625056, 840326822, 917498546, 751761984, 798449640, 1393540732, 1484933017},
    '{128, 1363946183, 2127733168, 1091187071, 722229624, 232690772, 2130043758, 868108689, 683601869, 1528784089, 629131781},
    '{161, 1649043291, 132870103, 101010727, 820887501, 1656774462, 560165759, 2061135611, 1518266190, 750000498, 1971492389},
    '{91, 396766448, 605905673, 157591805, 1845874584, 1006962417, 1593442498, 16332035, 838488814, 1414767558, 407852410},
    '{192, 17586756, 1197106914, 1196382383, 609065869, 1105993043, 389839119, 168737669, 927886875, 1929062138, 1032797798},
    '{132, 1407958825, 1347262099, 228549882, 239748890, 1920326078, 1569359469, 1835984585, 1600327871, 1882334368, 1020250939},
    '{38, 1070405349, 558491439, 2105103001, 912563207, 1027925247, 1795973433, 1402361302, 1888687010, 1810340124, 443954085},
    '{46, 1506101460, 1890282250, 785499655, 741668338, 1888910638, 498222835, 1041078057, 1269502296, 1613518849, 831572274},
    '{160, 1985008930, 1434354717, 1128740186, 892439105, 1043428601, 1854862667, 1634827717, 2014993538, 226164438, 1837293070},
    '{94, 1180716822, 2053182761, 601101282, 586925288, 104352683, 492407494, 1590331992, 110160733, 1931963999, 161604088},
    '{150, 1622313203, 1521447940, 238042234, 47793528, 988185383, 1625199102, 37138920, 75704342, 536941456, 233921705},
    '{236, 1041492992, 931974769, 676031667, 1628245146, 600390376, 1796274119, 4542659, 1790149290, 279038465, 1802799690},
    '{78, 1641645931, 43452579, 562818849, 479727368, 107773726, 72932823, 539953157, 829232586, 1072481097, 2015044807},
    '{192, 1684366902, 772414728, 1549082146, 1022807323, 2077291674, 1627353721, 410518840, 1315063390, 1376930537, 221215866},
    '{231, 235253296, 1774011698, 440553617, 364283724, 511559622, 470055653, 399640514, 1249689413, 1878195791, 506651040},
    '{208, 1796311371, 1142669697, 857639659, 424381106, 949975625, 1808561237, 1310780958, 237993796, 967274902, 1463978270},
    '{90, 1662586491, 531637849, 325997959, 1948182490, 834199637, 1322735029, 1432476818, 2028344898, 373284063, 1883901903},
    '{221, 1668118697, 2145210986, 4267837, 843070076, 6300876, 1107578723, 777368272, 1310335244, 1430598361, 1500743586},
    '{19, 852589076, 1041415936, 399977789, 1429283364, 1871443240, 246539231, 1463466804, 1722373214, 1942511973, 1617802048},
    '{68, 63101943, 1800854248, 1307789833, 1466653466, 350454610, 525351382, 1337313341, 1756514977, 1439271516, 1846401244},
    '{41, 1330839842, 24309825, 1715812580, 1055258368, 335898672, 1525356941, 462471375, 1741894281, 922781672, 1788281377},
    '{23, 1213269522, 663178661, 723482382, 761608918, 1033429485, 958948914, 597190258, 393873672, 461155379, 1777185632},
    '{119, 1037950284, 564241770, 1806350680, 504623999, 421137551, 1353923345, 1632379451, 1140057356, 768421094, 1467119046},
    '{109, 1321800146, 1718604402, 1392373970, 2012710511, 1096964094, 1116730874, 639516133, 559797100, 475403407, 108057831},
    '{197, 2036669414, 669567417, 1979422528, 457845495, 238089103, 333699074, 1868250881, 1088961584, 1939902492, 1531532782},
    '{36, 1643139914, 752603390, 442407373, 1513090166, 511690427, 217119515, 938019709, 2115555483, 1274304632, 1363774620},
    '{228, 1687611859, 1621892132, 2092155596, 1975523507, 794045607, 1317857524, 1555531794, 1884323709, 52951068, 1108911110},
    '{43, 1397263142, 1830676405, 2067220507, 154662993, 920045468, 135705930, 1593208847, 112179758, 1523898516, 2047424199},
    '{62, 24616523, 92815821, 1481274570, 1240799243, 304170380, 484309558, 657925369, 60615781, 177692981, 151128814},
    '{51, 1361297181, 303730217, 645183909, 858765232, 749634384, 485984505, 1081707123, 710844361, 1276908188, 664059879},
    '{235, 759000667, 1119997255, 2090874015, 778707553, 1217625520, 1587520684, 262678506, 98160839, 1446055130, 910770951},
    '{141, 1438779399, 722774537, 1466132623, 394699518, 1781787645, 1785588768, 2096400060, 1225729080, 1641400869, 1928907561},
    '{91, 1461698465, 451931501, 741507411, 275056913, 1644774869, 668241222, 613548422, 1929364582, 1183665236, 448039130},
    '{9, 361737349, 1153058658, 1591163713, 919830847, 420349022, 724864704, 1912744977, 1957097941, 1992260831, 1936679434},
    '{17, 1460871768, 1756573199, 809536722, 1984338552, 1091357071, 1338838006, 1505522415, 1817033003, 491588820, 94837790},
    '{39, 1960898376, 479026398, 1032237724, 1907969243, 381079919, 1711299326, 991249616, 1176824863, 1658775356, 118326326},
    '{125, 396091213, 1881399376, 1043664468, 1457991938, 1115244304, 319360770, 2115861263, 1599133044, 582007432, 2030582279},
    '{224, 1255724031, 955313073, 962432522, 767942619, 24743425, 1831024687, 290516910, 300904571, 15906485, 1687977804},
    '{123, 2022454266, 1388554513, 705206744, 1706585176, 97142874, 742497853, 1589832748, 1713429992, 1813861818, 1085319450},
    '{239, 441327871, 107547456, 1482941453, 951623633, 163684070, 463877643, 980166561, 709783280, 728921938, 237584135},
    '{97, 992793272, 310878491, 356990074, 1253060498, 1715557013, 1036510615, 145457484, 469670061, 1376530999, 2120573147},
    '{113, 149533028, 667177893, 978466912, 930708521, 1217631779, 1733071170, 1880799919, 298255603, 750272293, 737841124},
    '{44, 213021, 4375256, 194084620, 1114306025, 1150937667, 1475928260, 1081742459, 1321712366, 1833462890, 1730763945},
    '{147, 2034165010, 2122615708, 19515048, 1476716039, 1062936931, 619480678, 451718575, 1933574945, 1476309374, 1119610302},
    '{187, 213081097, 926490203, 684013107, 188896146, 601534723, 1824048202, 961451864, 2011045340, 1314122872, 234429869},
    '{98, 943740056, 1115913786, 1011835070, 1006165149, 54332088, 1113187148, 1755266344, 680736833, 487170459, 1556635205},
    '{154, 1700562593, 1582416228, 82173322, 883218067, 1541482554, 1334204901, 787368665, 1703440638, 504317164, 766895343},
    '{40, 799141670, 1118072487, 132812363, 1180848501, 1693945401, 597366080, 892794070, 1409132886, 1985299192, 387826627},
    '{209, 33129963, 1654992032, 69130063, 368254160, 441581135, 844764405, 1364802797, 2135627722, 681139939, 1174272721}
};

const rns_residue_t PTCT_ADDB__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{69, 1112177129, 533724018, 177369642, 1679005539, 53351151, 2070494231, 1541419757, 1696370584, 347098394, 437246425},
    '{132, 1073643523, 1839593152, 1737833869, 475564003, 1170319952, 1652591677, 1893033484, 1289139608, 1822810015, 901509049},
    '{57, 1573781463, 993476669, 1507418708, 874189345, 692173683, 1932035895, 102459850, 954571405, 326083750, 1858900645},
    '{129, 642013974, 330177291, 1879332416, 427739881, 26936754, 532533065, 238101500, 353341552, 1979250593, 1650878797},
    '{247, 1535568654, 1348127997, 1184988662, 775725998, 1284421050, 1875436924, 555592031, 1809645727, 421487266, 1836811102},
    '{39, 1805432572, 1479444956, 244255772, 1224792621, 319799473, 347843552, 36778632, 675486343, 2009285989, 294120590},
    '{160, 1986164299, 1598529120, 1436650053, 1643346751, 272751406, 2007774722, 709297180, 75598111, 559874537, 2069463409},
    '{247, 1573748398, 454327867, 1498198574, 2111692289, 49349787, 1863696371, 1862307614, 695707079, 1806252203, 285885356},
    '{240, 793712966, 1379276323, 940594248, 251432029, 1054277901, 1259679507, 1875681120, 94997645, 1179282860, 1651078168},
    '{46, 1175247393, 1859984809, 1570158002, 686201950, 1310180575, 224171677, 358778910, 1044836134, 1536609293, 996445963},
    '{256, 1209786133, 120134477, 542613025, 1303774553, 1945101820, 1838674287, 2099921014, 1995139141, 216989535, 1052103704},
    '{178, 323465262, 1919920335, 2120776926, 1636300435, 1539610204, 155259356, 1954766996, 585577789, 1447080485, 623930339},
    '{139, 1317357697, 563472139, 1848835297, 1030568413, 473560243, 303622603, 258042912, 1350930065, 1206935250, 2026007439},
    '{103, 273472673, 1009731303, 1449642611, 552032416, 1095771467, 1077074838, 2009540474, 1904124801, 1728187139, 39381265},
    '{13, 114973467, 1032654111, 424623647, 622386705, 958463838, 2083997397, 463044866, 1928399823, 1147380493, 1306913884},
    '{195, 205335063, 1886108379, 417507717, 1311297209, 1761787574, 733919295, 379871043, 1672289111, 2033261301, 470497663},
    '{247, 929474100, 931895368, 1135264551, 904652826, 26041372, 1282426129, 325859245, 285135056, 1076641535, 781758219},
    '{251, 2087640943, 111135999, 603708949, 1834610488, 1555370594, 2081115710, 1997540534, 1116957688, 41882368, 829777403},
    '{111, 1137914062, 1836344919, 520131276, 38364962, 1536109202, 1684360181, 905999782, 713215539, 474109680, 37534418},
    '{173, 50724856, 441216684, 1558450073, 175251215, 1427316833, 1325475737, 1883296117, 972722946, 591159604, 1257059940},
    '{10, 1790526298, 1142469265, 846814022, 1632341827, 686687227, 1030300000, 885556595, 300196477, 2118400296, 2120870940},
    '{132, 274699927, 251379310, 1526905371, 122336813, 341917247, 1485190404, 1444780683, 1826772566, 280136859, 99978012},
    '{142, 856480771, 1599804980, 2118686351, 2092037919, 747563729, 2060261768, 1561048654, 1061630523, 1455980166, 242505756},
    '{124, 1974415339, 119315054, 1564842321, 1660438747, 1550063704, 717930394, 1211259338, 1241714250, 793254046, 846536773},
    '{70, 143359175, 172540776, 932916070, 1922634533, 1868506359, 714680181, 1074790159, 1345953700, 2128692627, 202642547},
    '{201, 1117142210, 1679150616, 528529137, 1873055888, 2015238493, 718828362, 2144090113, 676470118, 96294373, 1772680642},
    '{61, 996309165, 1207918232, 807082959, 1936000263, 751961263, 1436729800, 1193790209, 2037821185, 1037098591, 1288545473},
    '{138, 833129397, 1902828235, 930672876, 228521519, 922443346, 1348733275, 2075808, 1161009866, 1292162685, 12766119},
    '{20, 790372, 81104610, 1539322725, 707502649, 575965510, 283699902, 347711999, 1982566773, 968607687, 205361198},
    '{89, 1697214270, 2070533899, 1249720437, 1338706745, 1732282582, 250645441, 2059198498, 566771232, 1647576203, 1653833294},
    '{75, 629085881, 617284009, 1259963447, 479018809, 57176881, 406981233, 299561556, 1919910668, 837949126, 392964044},
    '{66, 1155221626, 1115962719, 1107701070, 1884712944, 1906075554, 1485486613, 11167577, 1120042162, 567908486, 224547887},
    '{156, 1965386384, 269005161, 242053564, 610786302, 1838563798, 1476567249, 2059693533, 1777827796, 670852388, 844248888},
    '{2, 1134339825, 374409068, 1712228254, 1494014663, 1111161829, 111038965, 2002186539, 1207964587, 1283198887, 307022268},
    '{74, 951055157, 1324536092, 627027283, 1306671700, 464939953, 295729341, 828055863, 1213152908, 1335574469, 1376581909},
    '{189, 1540780196, 587249532, 685733135, 1621209726, 48171582, 141561841, 1252461035, 1787854826, 960780260, 1444163481},
    '{94, 1772712583, 82039703, 348823278, 1409838555, 1534338606, 1532893202, 536058282, 1312782605, 1973604921, 702817201},
    '{238, 684799168, 810617566, 1563868314, 2132277025, 1176205618, 1291617212, 1838737579, 1344807809, 205029332, 1054039331},
    '{193, 1957191823, 713610747, 1022258107, 137282310, 1747398000, 1678452136, 1374050502, 58494819, 1920146036, 1030312991},
    '{183, 1516519767, 153726826, 481122877, 1653785398, 1746494811, 1421695236, 1121160833, 1275308650, 1539636806, 333468000},
    '{152, 10127594, 1000689174, 313552564, 676065905, 622357239, 949605324, 384385279, 39249879, 1197981334, 949137540},
    '{194, 337931369, 1883587918, 2144223165, 855614651, 1520467346, 94829642, 1404149425, 1447443133, 1153651154, 1330699206},
    '{156, 2059688593, 1667457801, 1704998216, 212898688, 1283772960, 1816058199, 1838322636, 1715861534, 1275659244, 420883517},
    '{224, 100752787, 1003691475, 1891578874, 17834090, 760348900, 1518570040, 803557864, 289166598, 1465043885, 803412714},
    '{57, 1717345784, 1366360348, 23323035, 1158294019, 1463842811, 618382164, 2089062547, 323297971, 1548543634, 984931701},
    '{114, 937164559, 2051324299, 1359881548, 1048106072, 197283873, 1088081970, 600312125, 860429775, 1631863013, 873653663},
    '{140, 199733385, 1229119, 581351261, 400306788, 1275471543, 1314617845, 871309140, 507070491, 72930676, 264662275},
    '{152, 1535323094, 2110171527, 181617893, 1240107990, 1760785827, 625690953, 918847505, 1121377264, 913794679, 176667167},
    '{204, 1524898392, 328776342, 1478926205, 638627153, 1525155906, 190214825, 939014537, 1370006499, 1472770738, 1901673828},
    '{148, 1977356419, 1416042110, 1268940098, 1599005508, 1360518251, 1852933215, 1845618624, 1221987484, 1025654898, 2022986732},
    '{42, 1924168719, 1117521149, 1349322214, 1825385249, 722760803, 1514640851, 713033627, 1186258764, 2082051839, 665342042},
    '{194, 1624957882, 1323885445, 105666162, 1300983833, 1840544033, 1383379926, 922984325, 19271487, 270741065, 432310072},
    '{83, 1783258660, 1233720022, 2057058461, 932263646, 1711607144, 922882246, 2003002430, 1659266438, 1540243119, 1212675658},
    '{211, 767797460, 449130898, 487780479, 912922911, 805659668, 1076739181, 1976663147, 102864022, 1144022461, 570311395},
    '{126, 1787518897, 2129617489, 1795316463, 1508132779, 910772726, 823915451, 1567449857, 1749834906, 1936884195, 416712942},
    '{40, 1880538070, 1797055427, 1032899401, 28386578, 933519243, 2015643943, 587367817, 575599096, 963794549, 322785847},
    '{152, 1767143481, 1171034278, 801826112, 129903151, 1285551010, 98640459, 1499448647, 213863181, 990285516, 564816723},
    '{235, 349263378, 1725167867, 294977853, 1364875384, 1630016139, 20313273, 959416456, 1023240651, 844469708, 756943719},
    '{78, 287220864, 1433201783, 1598528648, 1239915840, 940797769, 922005843, 552867908, 180967113, 1437316834, 452718313},
    '{178, 1580529675, 230279239, 743086191, 532454816, 1607468248, 966242335, 501280583, 726033383, 915813203, 1232024914},
    '{92, 755984682, 825850527, 867645482, 741438072, 1015419087, 1868974263, 1280052164, 576935286, 1803245003, 862452203},
    '{204, 195958570, 1678176313, 1768673732, 377441428, 283910164, 714687245, 1414491619, 1114772996, 2038631762, 1235495759},
    '{113, 711514740, 1837214213, 1945467505, 605421544, 558182535, 716094237, 1114379824, 271557769, 2097514290, 1782698781},
    '{202, 707719628, 988967764, 2055368146, 1745192673, 177037800, 1835330505, 1017619763, 182878640, 546019738, 357572893}
};

const rns_residue_t PTCT_MULA__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{8, 1942190391, 1108279846, 1576746942, 1597202575, 1008218077, 1755696927, 26973342, 809216979, 758598977, 134595091},
    '{198, 27030712, 1512568157, 1594864172, 1111230086, 1818608650, 373734051, 1425137275, 949916480, 1269431672, 2087943425},
    '{28, 465477726, 504547342, 1194900005, 1241930234, 568467687, 758718919, 199048019, 161380257, 2015335251, 1821490389},
    '{41, 1412586922, 564032256, 268378975, 1495747516, 1274626795, 533485451, 1542347213, 1893771138, 1897328028, 1292225261},
    '{242, 436921533, 1483158813, 609360658, 1574599636, 2031732583, 384558370, 1232047807, 1425106467, 1930974176, 1705626134},
    '{227, 1528016567, 650615826, 278186915, 618307419, 1311308619, 548755814, 213782636, 922387831, 1898862520, 89279438},
    '{210, 583926293, 2081085140, 480937465, 1668466007, 147195209, 1987272133, 1014293251, 25123214, 558987147, 344777049},
    '{107, 1641468006, 670982100, 1529388824, 1622902827, 1494340022, 544883412, 2039038483, 1419140656, 1913065697, 701744729},
    '{239, 1959747509, 432237845, 2124884176, 315055569, 1699063430, 731896631, 193975114, 132734519, 1394879121, 2020923004},
    '{32, 1463714210, 370675717, 1083624262, 2063233576, 159758928, 802007501, 1049374078, 1500079406, 866955350, 1322825414},
    '{52, 513250233, 1682219412, 285973292, 2134541180, 1884162796, 1890500604, 38510875, 688505642, 191329257, 814282102},
    '{180, 1061319129, 783258884, 1808230938, 778146593, 1940754352, 611117401, 1332512294, 488229555, 724640537, 1036597523},
    '{88, 2114792783, 770884458, 388457775, 700688312, 1832745982, 1948302522, 1614386281, 929619194, 2117016003, 769431272},
    '{72, 1012456776, 1583622373, 875020987, 1667911781, 657628851, 711575692, 1303143889, 1129611235, 348798143, 1889933972},
    '{133, 1004221052, 1709247619, 1427389829, 22920052, 2106634293, 1533207278, 450021336, 770097250, 677811438, 1092521533},
    '{210, 70553642, 1400778590, 951946558, 2062486213, 1103658055, 471665880, 1403476042, 1010497471, 67984491, 2112839143},
    '{132, 1001671948, 445786164, 506704613, 1716568504, 1299289311, 955263382, 1595769511, 2044946777, 1703692673, 1180399372},
    '{18, 1232095861, 749614638, 1830863092, 2036390604, 1156789167, 1456057091, 406015008, 1416964753, 1677230307, 1369258496},
    '{22, 1850328528, 1370702567, 1005043130, 872891855, 1686880939, 1587224344, 1547268841, 921038592, 606025281, 846262707},
    '{176, 463010642, 2010557684, 1838551958, 1042119197, 2074131871, 2060070898, 1731875445, 1981261671, 528674814, 1876818729},
    '{106, 760105115, 403335344, 57467873, 841283704, 1289474371, 1157999700, 382366238, 1378319343, 734547338, 288595126},
    '{54, 1627103418, 987875026, 464686871, 428148530, 1843410813, 1892019922, 2010067432, 1113566974, 792514675, 1441199601},
    '{96, 1644661273, 1111461232, 408374328, 1921360797, 821748707, 1893640589, 5381847, 2130104734, 731473146, 53720790},
    '{57, 1345103202, 1123560672, 1550172287, 832190747, 223261778, 139373251, 2133910276, 1835094491, 1932005028, 2002590692},
    '{210, 512896762, 1102785639, 1706891565, 1023585571, 1419279740, 778712040, 709917936, 1114620877, 1610698132, 32401113},
    '{203, 470826664, 125927288, 2079166366, 1058774623, 569171239, 126748747, 1157759190, 1995028150, 921135910, 955692235},
    '{240, 679342269, 1874053283, 689022283, 1004653433, 874393063, 321273502, 907792174, 1453914479, 1882187540, 530389187},
    '{8, 463044738, 686131157, 1171758372, 912781198, 435791355, 1263560521, 655021659, 924866292, 959961362, 273626562},
    '{116, 971086429, 502824611, 1214101200, 377507706, 2124496024, 91067571, 1849699526, 1688093211, 513641623, 74525429},
    '{31, 2053403198, 492340494, 1594806078, 560014570, 1501298268, 1127783486, 1465766363, 555644378, 1393572054, 690444514},
    '{225, 226561171, 1149855034, 512094522, 721790648, 1088969298, 1389509648, 631510851, 1259066450, 1734109602, 1144570067},
    '{165, 1570252194, 2097200994, 1692094388, 1450194159, 406521305, 1744081060, 483101481, 9221368, 123186499, 1227588526},
    '{214, 1245576533, 951461981, 1555536358, 22455131, 1160036085, 1229733652, 77572072, 1580930473, 1507791573, 1202801219},
    '{121, 341483963, 1353277146, 1644304409, 1260005987, 1147626585, 1504800720, 1278044279, 171439070, 599330283, 1047288078},
    '{157, 935858047, 328852992, 1543979028, 829829116, 316139328, 182328946, 1557112417, 930755190, 1420953924, 455841514},
    '{69, 1097473864, 716529564, 1477123785, 909496980, 1477285728, 1360389893, 1068730160, 2142488217, 69898309, 562662700},
    '{248, 1151822374, 892779787, 436778706, 550903815, 631572305, 1248351819, 1659941978, 1391141631, 1466561210, 2003192767},
    '{11, 855184120, 1370594143, 450011415, 259170187, 1999540980, 384904475, 1061641772, 61847415, 547684988, 1465225758},
    '{155, 1510507786, 2034614154, 273043917, 565474730, 1669062975, 2138482399, 1922001852, 232526906, 1652759080, 1017452812},
    '{93, 1925585863, 19459817, 1682091932, 1552118739, 318392172, 192506187, 1940435872, 123438689, 1328858365, 1256090260},
    '{54, 1902488394, 1785541943, 1133281581, 1282371507, 2025281498, 1547942709, 255577034, 750446157, 567005069, 398301184},
    '{67, 23399313, 466590924, 757630496, 1022805572, 1341235758, 1466124152, 1323662442, 1766108061, 174336621, 1010990210},
    '{253, 1430670404, 311478755, 567996785, 1052786410, 1379130681, 1845845794, 71436116, 958705728, 956605410, 1338599945},
    '{198, 1390710378, 1037570678, 1108904473, 1677741669, 857662708, 350398909, 1627359010, 1503937793, 138184202, 1169090343},
    '{31, 201656612, 1286451214, 848042304, 776074879, 1399714152, 2125884377, 575104360, 59239751, 1560416545, 1637058886},
    '{251, 927361747, 1701718228, 1795242901, 1779477708, 1412719922, 1054743111, 1632221061, 564594104, 937011291, 876219167},
    '{223, 1847833898, 590073939, 827127171, 1889519548, 1313453354, 726193472, 222568959, 423413860, 1985065105, 367486078},
    '{69, 529017193, 900096154, 740699088, 249636548, 844701223, 706960671, 779395157, 1795225449, 309716365, 70431762},
    '{134, 1958995591, 1310974804, 882813132, 214940834, 184262013, 1976288674, 1835991750, 835295653, 2064395812, 1651972558},
    '{56, 996274519, 1290181822, 989917541, 1930073436, 115362574, 1537368246, 635377968, 1471930933, 522823383, 1247365939},
    '{16, 576490156, 512285100, 1945163198, 917209143, 565376799, 1553405500, 1061772778, 1764499394, 92616979, 1895811105},
    '{98, 849390055, 1379771065, 633360087, 1001451787, 736810443, 20479084, 12231279, 1801451460, 1361276559, 987309191},
    '{25, 969541868, 1127432565, 1009577519, 1250205410, 430983820, 2070418361, 801942769, 1746560923, 112652101, 1815872312},
    '{133, 1496887334, 1787761355, 1661172363, 87161841, 1166800670, 176968537, 313641114, 315872045, 1855369291, 1726860247},
    '{255, 707317899, 1716445887, 498899653, 397367423, 759963217, 377257667, 232152487, 1523597715, 294285404, 1246726735},
    '{209, 1753290389, 2110929985, 342956106, 362209076, 437600733, 1371149371, 1758933564, 907806461, 1240467885, 715534427},
    '{137, 533645219, 568786819, 559535281, 787465107, 1443994323, 1455814553, 2135398214, 234380350, 181222162, 304332736},
    '{248, 1394927139, 1852530546, 1083179886, 964068144, 1402411020, 810746584, 920422169, 781928358, 1363047124, 131740875},
    '{209, 1509014639, 2090330215, 775465805, 1986136158, 541493795, 985928363, 642653347, 1994499937, 1935728719, 961443594},
    '{84, 451027032, 2020571432, 118724509, 1144152806, 854404320, 537383627, 1179882939, 1207828566, 839251482, 1587041376},
    '{205, 1149362546, 1419674770, 570539415, 2118653666, 480062570, 1596938904, 1139219480, 462159707, 1963550289, 759871044},
    '{123, 385159668, 1801525800, 41192683, 934778930, 44989731, 834305578, 925913700, 1516050815, 1168697275, 980707067},
    '{185, 1104134728, 2046171241, 109778488, 1788497180, 1331328145, 1157729574, 28938652, 759808047, 844739977, 879013258},
    '{101, 724793418, 1265830116, 338075706, 894218798, 193179462, 1552331807, 22014586, 510113616, 1490660771, 1857905391}
};

const rns_residue_t PTCT_MULB__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{174, 134237389, 1428005063, 1097395299, 1032973319, 1621760884, 566734468, 1494808512, 740809603, 128054418, 1044818298},
    '{47, 1343530766, 1368748219, 1270271977, 1583322503, 716763227, 670830818, 126615209, 637328160, 998160139, 391668259},
    '{188, 816702889, 1319256226, 1613152897, 352164695, 1677602955, 138114953, 645934063, 290395768, 839098413, 764451793},
    '{226, 283068568, 1739728747, 1127694320, 2115436676, 1952733916, 857382157, 453960536, 71177508, 631468363, 433659745},
    '{86, 2074653264, 2118038288, 323469497, 670666572, 854303481, 731755072, 1421533891, 1220061146, 328940405, 696469293},
    '{138, 317896598, 2105503523, 554584923, 1979863592, 1400276934, 1547255884, 1629588531, 985314321, 1326731271, 1946713594},
    '{252, 1995677625, 278638278, 1912012264, 1631396399, 1412445072, 1489113591, 1178499611, 1129785115, 1045281546, 565962545},
    '{19, 921222581, 894082956, 1133352666, 359149632, 97799197, 1824988679, 987464762, 1445469841, 680201948, 711503236},
    '{156, 1858778257, 1139579280, 289920282, 1006110217, 1702290610, 1076724870, 1443189408, 1099464161, 47426085, 2057179475},
    '{245, 1612197821, 1881980401, 1970182752, 563940917, 2017017273, 195316922, 1744448243, 1843709737, 459485690, 181153704},
    '{105, 1637356508, 949865368, 743380049, 1829304193, 560203748, 1723981730, 1139651097, 1035304402, 969845664, 437048446},
    '{2, 935933070, 396929573, 1529671135, 659746486, 1858298434, 1546688379, 942866216, 2005857427, 1024825256, 1930671610},
    '{200, 1523825169, 1167361788, 171767121, 822014966, 213164029, 1378074615, 1517793717, 368188988, 1626427128, 643171831},
    '{117, 588348566, 982732225, 1211890992, 1178942455, 1305735229, 2041824115, 274843865, 1240774053, 1831307258, 1108447262},
    '{171, 1324152047, 1939021540, 674008712, 1729916942, 679117970, 1368762257, 1947602191, 316390891, 2040282209, 6779823},
    '{52, 1287363716, 490273852, 750744871, 1622982767, 735731509, 2086866443, 1314683198, 2119252033, 658227941, 169487950},
    '{92, 1577176414, 1968967151, 599226609, 1027723801, 1396080577, 1587803278, 849992874, 731646952, 786495262, 1215467403},
    '{236, 1047619584, 1968365796, 53588433, 1620368998, 379356405, 1448830804, 1589774942, 1092365228, 810662780, 1027167485},
    '{216, 1612259907, 1161841172, 1955708606, 1709776988, 912771389, 1239980474, 1847505453, 1104294185, 1835520101, 2101113129},
    '{19, 1743802230, 358201882, 2053273982, 1434287024, 1598907671, 720282067, 108893791, 1637814715, 739616652, 1214303061},
    '{231, 157861518, 1853653290, 542162241, 1027265338, 485465462, 368367381, 481446590, 1770055702, 1998165999, 279954230},
    '{142, 1253117584, 1612176876, 1486122682, 913049380, 1846245480, 937420488, 1001816750, 529981300, 407125185, 571524193},
    '{68, 628574548, 249619774, 511728562, 1592551111, 1523286734, 885353279, 1708532610, 688156689, 698108794, 548067015},
    '{84, 1172264309, 1203877326, 715038614, 400755224, 1623074631, 1145858594, 2091942845, 1096624147, 1701039000, 696730846},
    '{13, 259316138, 826108446, 1797289825, 1562338303, 451596947, 1023383062, 1521750533, 1409717351, 1167585826, 2070557107},
    '{188, 824230468, 1704303499, 1751134133, 2046951024, 278374459, 365483332, 948392678, 999027232, 1513202181, 2082486656},
    '{252, 1308844218, 1218007083, 794845621, 993427253, 1837906142, 426095872, 2105779385, 757080333, 895788425, 2027096592},
    '{66, 134614386, 504048122, 1306513325, 513461409, 2050499918, 734145528, 953837837, 883887465, 429361258, 1264943985},
    '{172, 531730472, 1465712037, 2746989, 240099497, 38066992, 901974107, 1128472243, 971893001, 1977971285, 1470187373},
    '{183, 348156718, 292213124, 785757356, 1218424772, 1066994678, 1303375060, 1897333919, 953131564, 1397261904, 1399318585},
    '{153, 2091762075, 1692416176, 773644586, 977626107, 230515669, 1051590281, 1980698005, 542109655, 2041444373, 337196556},
    '{205, 894467761, 1027563456, 1281598520, 370239477, 2050792549, 1696367096, 2100753701, 1762017500, 935053612, 533379783},
    '{100, 1655207864, 290628874, 429408233, 1617543062, 1679508465, 821517053, 600233808, 246868592, 731241919, 1458474433},
    '{106, 1103063546, 2050746808, 946783625, 2084599031, 2049776500, 247439523, 969342383, 1450199214, 1311805298, 332643696},
    '{22, 1833693632, 866604638, 2132268812, 313837518, 653078579, 100104031, 434843436, 614721496, 568446582, 1114570544},
    '{154, 1554895796, 341111030, 1049774995, 1592825892, 1056679059, 758402742, 1102929241, 944804941, 1820413985, 21354376},
    '{208, 1159778120, 1576002010, 613322685, 2084384404, 1787495918, 1426215631, 2036989877, 948970666, 1134078720, 125888604},
    '{56, 1885200337, 2117816217, 188057812, 705637282, 1168141000, 1307204226, 519746529, 1780278795, 88477105, 957218813},
    '{222, 1025951530, 428914736, 1898618019, 143512564, 1259923531, 1028234748, 1150143168, 957312947, 1193085676, 1086537222},
    '{138, 1953450941, 169623642, 1666676572, 719564066, 1793128865, 367242566, 351773842, 351610077, 1676925950, 1547117518},
    '{107, 195477158, 1429983969, 840324779, 1748647681, 26184609, 682120763, 599738788, 1551872442, 755002740, 251342226},
    '{7, 1189050730, 944458208, 900511868, 222549191, 752414222, 421418882, 1869847280, 1864898375, 98898434, 1575062899},
    '{217, 2121886737, 1322754944, 514754965, 2012182906, 393300914, 1606557611, 1353236568, 1297064395, 2137767866, 1652109812},
    '{22, 977102035, 1645384411, 214723943, 331977999, 922424158, 1457203221, 1383407936, 596798105, 408458523, 1609270183},
    '{29, 704160994, 1270310833, 1081449351, 1482824079, 1820667023, 107749317, 552971288, 1324619273, 192625045, 279264417},
    '{215, 840879971, 70474609, 1194520857, 387140281, 1721165250, 248667599, 601303381, 989146752, 549538435, 1708846752},
    '{61, 1056581703, 497414372, 1647980591, 1354572418, 47990165, 1613646486, 295037373, 1246972677, 1426056251, 347984294},
    '{34, 1270965856, 547530648, 293426884, 2055150284, 586811133, 2017396859, 1776837448, 1959852432, 1300748659, 1255701836},
    '{117, 1788457010, 654374293, 939648935, 1222681673, 1654064529, 339944985, 1340803943, 2124346521, 53153255, 2059131892},
    '{88, 426184100, 724040560, 1551703035, 860956391, 1334518706, 1111372456, 303984095, 583323394, 1958138183, 1406477208},
    '{233, 227982169, 579774783, 1841482286, 189866890, 905497901, 1883877768, 1266337621, 1119118896, 1316477123, 480828296},
    '{92, 602345686, 1613299457, 412524636, 228456342, 828754188, 1808906976, 1091549077, 1576732961, 322512709, 634581523},
    '{254, 418392881, 796004915, 546131794, 2119730953, 1920476884, 131308055, 423886527, 1185437003, 421506085, 137036434},
    '{170, 1037791958, 713394074, 553187872, 818243747, 1634333509, 657444721, 749376026, 528301747, 1352515263, 1654459218},
    '{37, 509937076, 735213544, 903128474, 1963205359, 506646608, 846337614, 1339912611, 357409041, 1668868310, 74627100},
    '{111, 652325240, 1563614897, 1933504357, 1767610416, 217514640, 478923985, 1260921035, 297454705, 1363194724, 894244722},
    '{137, 1965202222, 415611235, 465769792, 1004498435, 1333683169, 380667588, 455716144, 2140867716, 616453975, 311720381},
    '{88, 1704933659, 471248388, 705777320, 234350856, 493027799, 1880715131, 347176734, 243284979, 202539139, 1248962491},
    '{150, 1803446067, 531228489, 885945778, 836696200, 460856497, 780636889, 253609912, 1886842558, 598705405, 1374611672},
    '{81, 486331132, 259442841, 1244558980, 840568959, 433391025, 1526555807, 1796925910, 1325146170, 1474418563, 198217415},
    '{13, 91212659, 160312205, 320291470, 888293732, 1207411456, 982148156, 122083268, 1706414990, 1363924421, 907533873},
    '{122, 386533143, 882024002, 1434226632, 1387292814, 869874323, 200007975, 2042048837, 1696841881, 625486992, 1851338223},
    '{243, 921031490, 1726284915, 2134692199, 1161652340, 2009676127, 635600466, 663168876, 1725804627, 401218360, 1137007739},
    '{22, 671443214, 1585783215, 1850580188, 1889677642, 105606530, 1362831329, 2004099051, 1137214276, 1793730808, 409151585}
};

const rns_residue_t CTCT_MULA__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{110, 1299346805, 1403782299, 587003490, 137848143, 563378774, 1148054741, 1195290417, 1746578989, 923920916, 1994815838},
    '{237, 419002243, 831183066, 714331155, 461771381, 145902692, 876276914, 408015013, 1828773577, 989851997, 513775740},
    '{118, 218118354, 1019622526, 433406246, 76447640, 1508232887, 2019092901, 1807367968, 922113072, 1539668403, 2095160406},
    '{192, 815928782, 406691916, 1842173433, 1158409485, 933531943, 217381044, 860465039, 1793627267, 1496062076, 518178337},
    '{3, 602407404, 836561216, 1837820231, 861392792, 536863546, 1906139361, 939821615, 1574746174, 445189491, 955174014},
    '{38, 1942004599, 1248662899, 331669436, 1771043321, 1076769762, 532990289, 1889646424, 1549366017, 1327738856, 954818080},
    '{121, 2090889630, 66190353, 1494597117, 1412911675, 568936137, 1783910778, 2015318647, 1305260790, 794807879, 1975341860},
    '{38, 806279690, 763969110, 1638687697, 1650890823, 598088115, 1891900701, 1437849668, 1185730632, 2029394491, 344451105},
    '{59, 187779813, 1992696656, 1969894273, 245513665, 1792926493, 1731702788, 1834686870, 1604528689, 544618900, 1541008745},
    '{126, 2035466254, 231232247, 1291181876, 1755304355, 1244063041, 344977647, 1989741272, 1171997083, 1453622684, 1812274778},
    '{221, 121109328, 405422839, 621567688, 1013424413, 2099910405, 1262750558, 890943996, 1449683297, 1927040586, 653408876},
    '{141, 1617653448, 1119475365, 560153801, 1710786672, 452099244, 1425767102, 1247613295, 816463989, 580373801, 596759735},
    '{33, 353559758, 92128392, 719540503, 1355776254, 2013269200, 1352222026, 1787626865, 1506984291, 1206481344, 1515825621},
    '{148, 1869695799, 1665387801, 43864939, 202899798, 48510580, 1616139006, 1246613506, 1102624837, 1802042495, 541314464},
    '{55, 1402611723, 287036613, 1848819089, 1450978882, 904270800, 1537022645, 675879517, 230173479, 928835985, 283659236},
    '{136, 401536998, 1075346043, 1927610629, 272409979, 132860498, 837072811, 1234841185, 1050244356, 214993005, 1528206370},
    '{24, 1021098566, 2008740718, 282667552, 309390186, 46372921, 176079607, 435105446, 882879309, 680257662, 1044729788},
    '{85, 1180037206, 1116541672, 1026104252, 1373134753, 366032232, 46643658, 66333895, 1194899753, 963855510, 1877883232},
    '{175, 447805553, 190154466, 1162248893, 172170252, 1292590917, 1124688666, 790573369, 1233692802, 974402479, 1787136199},
    '{72, 2058938150, 1938046301, 702121852, 1737707815, 872094299, 1638198367, 587023349, 803263155, 2056812401, 649343668},
    '{146, 1236633399, 1267428485, 492172553, 817775714, 206666521, 934978006, 448041759, 1544893342, 1352581606, 722275096},
    '{203, 1239699069, 1874812178, 1231551617, 1749155321, 141550309, 2035074916, 798627633, 1346275158, 269516652, 392588417},
    '{146, 101060542, 702049416, 54423482, 528938447, 1692367388, 1899516935, 156516640, 378366033, 1065629079, 231321712},
    '{104, 2061582806, 251784306, 1377208939, 158840716, 1496901061, 800093215, 1466500852, 998861769, 1112691879, 1293287902},
    '{222, 398801077, 353047515, 1851281786, 2135720201, 511175065, 1336887217, 24343392, 1678738147, 1788193454, 313870142},
    '{104, 280555922, 2041580318, 1930478057, 584190896, 1771108277, 1387273587, 161470239, 1312213928, 1809157344, 1495501978},
    '{209, 1577953301, 1698613367, 1451986886, 1251467187, 632114648, 1804371031, 602999691, 463556136, 1566488337, 1592099534},
    '{107, 1911729906, 2144257412, 453983101, 1347253978, 1408788050, 1276882461, 1679871305, 1285131764, 476664029, 1053342306},
    '{128, 2079192547, 1355369537, 1046847099, 704299639, 2008435448, 1637072275, 1328422346, 2100452359, 419231915, 371850414},
    '{45, 1046764072, 635823394, 1254868730, 779608299, 960061927, 1451629425, 1220457344, 684574526, 1704729198, 1436344271},
    '{85, 310479079, 756331814, 396691956, 1399199049, 1593242608, 1664942870, 1714026399, 1697194997, 829836092, 544965237},
    '{199, 1869053282, 2077572138, 1141757943, 1632619954, 456284670, 982914156, 1031923441, 920750754, 832630167, 1043339379},
    '{200, 1455920191, 637363102, 902886411, 1320758481, 542562838, 1469730718, 2061424076, 871172886, 2065645201, 1918286142},
    '{87, 107213630, 19435748, 446659178, 1043103882, 1861795831, 563413998, 1658061775, 745080054, 937049685, 915763200},
    '{154, 1578461463, 120368646, 2125628132, 717666189, 1873637731, 1677191171, 117784506, 507245753, 852279113, 1686708729},
    '{221, 1356996973, 280556542, 1235240253, 1460918527, 658047045, 364307078, 781146195, 127276327, 618755103, 149575259},
    '{44, 248290576, 1062504122, 441504959, 702277791, 1001769440, 643403661, 1889151793, 81092274, 584998935, 1649053086},
    '{96, 2039822495, 420187232, 1350887691, 237004029, 315466740, 414881718, 1185931239, 1236670628, 1574739309, 173540443},
    '{178, 1012628469, 342176616, 2026767076, 79959364, 514993075, 729549499, 812807307, 608335849, 1851376932, 324629726},
    '{122, 243164514, 1612919858, 1159323032, 386420383, 1138862644, 749619430, 935675839, 1243223812, 713279809, 397461180},
    '{51, 271114718, 1599516531, 445557031, 769437225, 1900696335, 596165543, 759652897, 152759070, 1301385492, 1041995074},
    '{28, 144471336, 351091548, 1541847922, 614489496, 610844737, 1653195252, 251521464, 1189812204, 567960843, 4581957},
    '{94, 1368231850, 350982889, 387380442, 1660119531, 723829080, 249658364, 1712184500, 1613380748, 1294139270, 1485963651},
    '{206, 1653541345, 1793319285, 962980114, 1180695586, 767709351, 1755153684, 2059428819, 431959771, 1705355775, 4785818},
    '{164, 314115718, 2051266120, 700117885, 477611727, 2098890655, 1555049784, 145987970, 186138321, 66178701, 149897604},
    '{232, 1981345765, 110182736, 2037526135, 905884912, 878190374, 659077779, 1123312379, 605627621, 1800950368, 970963232},
    '{55, 1949812790, 1122740616, 2053242190, 1744005388, 92715243, 1967528710, 456008743, 1688149928, 1639009864, 2132085569},
    '{79, 70015732, 993954977, 1633551774, 595208967, 1084547173, 813127300, 1189562117, 734563850, 1669244455, 869686648},
    '{148, 826171215, 905953770, 1178694995, 710854743, 91828568, 1386267235, 2066307411, 1433618427, 908639041, 1549106943},
    '{154, 1690694065, 48096440, 848885011, 194378449, 941878882, 2124878488, 1626075184, 1583650054, 1540152306, 962507813},
    '{152, 593141016, 1596585315, 1429648758, 1021605114, 1848222131, 798657859, 873278854, 1472603605, 2027558394, 915553169},
    '{146, 1725294593, 640352198, 118835163, 802803531, 19029412, 239825698, 132597629, 2059638412, 733348652, 586411465},
    '{192, 1022090647, 1546172643, 1718787610, 1919002022, 2037968170, 492865805, 431698590, 2002513365, 604625649, 884073435},
    '{189, 1143800630, 1554925210, 718459140, 1667254507, 905902665, 1587011375, 1592154242, 1890469638, 1976197398, 1498493846},
    '{94, 1944064900, 675991317, 746839625, 793128640, 1667366775, 1421083199, 359630711, 484915829, 345790357, 215297993},
    '{5, 1654360801, 1023788744, 2000720166, 2052176393, 1697686366, 168850960, 850582077, 2090351704, 1738410734, 798274497},
    '{119, 764124293, 56639793, 396350036, 1988320671, 1754080874, 500246174, 713177001, 376787754, 802264962, 1151776831},
    '{22, 5463274, 1396871004, 15294220, 1021127834, 422749043, 2102448275, 1158271956, 119806902, 639132385, 143660195},
    '{29, 403992134, 642688285, 1839944497, 674572373, 131127082, 1297715504, 1379292174, 1288161079, 264729622, 93578372},
    '{16, 420775520, 455394450, 995878876, 909619465, 1136342543, 1335199267, 2030257217, 1182870568, 1180584879, 722251706},
    '{202, 2136181068, 1007091116, 1060242500, 355433225, 168190043, 682726543, 283923484, 638866985, 1429163714, 2023717914},
    '{193, 811240577, 2095315097, 1697121281, 1655254286, 79103867, 2046434274, 705824547, 1724965403, 1027886396, 1858305364},
    '{93, 1322934947, 1746316738, 646826661, 1591374453, 1594918446, 1570576224, 569834171, 154207366, 1491479512, 672900208},
    '{10, 1150681445, 842425171, 142143331, 1694490784, 690933188, 620263165, 104490636, 605682000, 1300742407, 907837}
};

const rns_residue_t CTCT_MULB__GOLDRES [`N_SLOTS][`q_BASIS_LEN] = '{
    '{230, 19934924, 203821313, 1794224652, 1604800850, 1763858360, 1460600622, 143463322, 942294528, 1017362565, 448966085},
    '{158, 524066176, 361939837, 1574111696, 864517083, 212122131, 960909550, 1706985495, 285228610, 1750541756, 754013373},
    '{0, 1197390161, 1602243054, 1466136873, 1970082760, 2097257266, 534757734, 258599115, 953097602, 51007536, 972345865},
    '{18, 1582256627, 360916998, 1398866012, 298004288, 551047351, 35534951, 165334963, 823039020, 1553949158, 796571965},
    '{61, 1645324975, 791426283, 439002269, 541363314, 141592247, 666696878, 214469798, 1486686286, 1019147306, 1751164870},
    '{240, 1599668221, 1472635279, 480264335, 2140383729, 624343888, 974165116, 1088219441, 384968604, 1101105177, 311696121},
    '{133, 299705862, 594156348, 730263544, 50114150, 1417305244, 658640255, 636040295, 1003920527, 117871298, 75642625},
    '{95, 676233315, 1919398033, 1383029022, 1435558568, 616440162, 609631632, 1874937817, 619268211, 1725973592, 1201769942},
    '{129, 652396528, 275865075, 1231418979, 1703532142, 235391250, 592097874, 779268367, 361532710, 811545851, 1436530877},
    '{40, 236913049, 636417988, 1221376810, 132522850, 581666584, 1960167916, 221910010, 1684031467, 1771210536, 1808748134},
    '{58, 228422679, 1526984371, 722919429, 2144094048, 788805229, 1510755809, 438254285, 15678218, 206236511, 901984165},
    '{140, 312722292, 2080437056, 767627814, 1716936759, 1017335470, 1073939605, 1635520461, 1422634208, 1051426187, 1572024695},
    '{198, 2146235373, 374410586, 1173256091, 1271382710, 865461045, 1484720209, 1961905024, 191528816, 986836565, 1483604290},
    '{105, 1781087047, 1133058910, 662837221, 298116656, 2064542234, 1470235807, 1665099816, 889345969, 1974351645, 803261675},
    '{126, 1216183406, 199681306, 1341319039, 1070621072, 393653416, 1873077417, 1027049833, 2079456823, 1582700386, 698036157},
    '{2, 1192984654, 1102440738, 1286074067, 77637294, 50940435, 1609611341, 895655626, 1169858575, 1781567159, 322035543},
    '{46, 2114922228, 983564552, 1890461788, 1865698893, 906975301, 1950421792, 954526427, 227691145, 820733688, 111905522},
    '{170, 378063470, 1989954905, 1334406903, 646796025, 152180150, 614060403, 1591333982, 956620190, 8312255, 2025745096},
    '{11, 118113708, 611624453, 29842820, 1346022494, 1832938598, 1165383781, 763242191, 1460088355, 1399378753, 2030744455},
    '{78, 147022588, 494427424, 529718654, 1295312385, 522561525, 627666286, 1762714530, 831111675, 824949267, 1365367804},
    '{102, 812871209, 1798328280, 1453486425, 706974145, 368056581, 1150054668, 1025337181, 1729291294, 2049915648, 1041313109},
    '{151, 1930832964, 506320116, 1439655418, 1420488324, 1966357347, 418461866, 1356108325, 338064760, 1138356998, 687986101},
    '{66, 1457933953, 658203937, 589792889, 907387054, 1670266715, 1239988934, 44282732, 772055921, 1539947260, 1851817941},
    '{59, 818048509, 1639532431, 1806315367, 749706519, 874634001, 662214784, 665567255, 102269774, 225856375, 230889667},
    '{73, 1465654507, 1878805961, 948935012, 1826410335, 1815394594, 2018867854, 798960790, 1235008674, 1981007187, 153854679},
    '{76, 1982009497, 726146221, 1876035951, 1926244322, 85148385, 815716686, 688321467, 329792215, 967352960, 1434128236},
    '{3, 337915003, 1686581354, 723698839, 585761487, 1901134876, 1747853779, 740656829, 883925456, 1887039315, 721837912},
    '{254, 1289390678, 1648102692, 547670781, 492620967, 2014201916, 1287352404, 1088061537, 1086362838, 1766364293, 421348516},
    '{74, 248665296, 457972021, 1867624259, 206071637, 66272155, 2077945086, 1456015323, 836214734, 1819670928, 544213265},
    '{186, 881038927, 365216635, 1568785574, 455218157, 1063346420, 1211486860, 1706842226, 2087172485, 928891656, 479573231},
    '{126, 2054899700, 626679175, 834020435, 1276758735, 1705445499, 229411077, 1760313484, 78380804, 943253661, 1818964014},
    '{159, 1454532051, 2015452537, 1256674454, 398714238, 1592157178, 1315464039, 745423128, 2544072, 1925099198, 1160014698},
    '{118, 2022647573, 1157271137, 976845443, 37273486, 453990176, 1794367146, 502750189, 1045722364, 220384919, 2137799129},
    '{110, 1438298075, 503037433, 1972956830, 1607371024, 1889515483, 974881099, 1564278768, 1092315393, 1694070264, 837669016},
    '{87, 1400889797, 177792067, 1065778747, 416114075, 1234969352, 1283978880, 255724309, 1452910240, 62247110, 535391687},
    '{195, 397653870, 1131019264, 791912879, 134510158, 21650119, 212600880, 762847192, 235213277, 883654329, 1042142706},
    '{232, 239404217, 1487886224, 833713396, 1621289470, 2144336776, 1618489713, 1725999126, 2088001564, 944985277, 841903732},
    '{120, 1837166903, 67082533, 1304211787, 2040864169, 1272791810, 787802443, 2146904905, 1169475022, 1919227674, 2010890603},
    '{248, 2023363861, 1143292110, 1814598857, 724748061, 1756062873, 871252556, 1397073569, 384397517, 375270723, 181042463},
    '{136, 1741535254, 1704003775, 1251917991, 1604368174, 1507946264, 1540622299, 1092905553, 392789421, 1688294536, 1298619962},
    '{33, 1673796651, 965440144, 1547419035, 169194326, 383643572, 1830864628, 602455932, 322493846, 1182972478, 1249442749},
    '{25, 1315328258, 600274022, 763157781, 1650818294, 934839164, 1116802720, 986898392, 1072707820, 578555610, 174389582},
    '{26, 3316726, 1290633603, 1951611536, 53311718, 223405178, 1074929908, 358157200, 1826567113, 2033966666, 1787244981},
    '{139, 416605210, 1009793847, 760490556, 1967503237, 400331693, 1112108412, 998814841, 439396702, 1164817130, 992483776},
    '{203, 471340415, 1403328240, 1114720737, 65042372, 1836101608, 1980344127, 1176540714, 382738590, 1163271949, 1189442645},
    '{210, 1876470598, 2100592105, 1747883308, 1104174446, 1554621658, 1491092218, 599872700, 1616842804, 497611062, 1188931380},
    '{73, 1843179803, 934403001, 958919574, 1075331317, 768941419, 552652423, 2133430879, 1210419988, 1936557000, 1962744308},
    '{17, 1879923187, 289239480, 991003781, 571736878, 296209307, 458437606, 989036081, 2118339765, 1218974240, 1620113896},
    '{130, 1875660125, 80412405, 1163845320, 593505254, 1882560135, 562820228, 607143779, 781676795, 760592859, 283669864},
    '{256, 1418183370, 1984828179, 1953120276, 831709750, 1863740799, 202574356, 1776480790, 596741165, 346747878, 25705924},
    '{54, 1983645311, 1247325447, 1056160302, 892164020, 625497961, 1436515195, 837355041, 17542047, 2065075189, 706212235},
    '{64, 498498184, 185146808, 1361083023, 2017756579, 404077717, 279728516, 1295305092, 250367439, 1432656235, 1051475101},
    '{109, 1819312988, 1370619907, 12603677, 15537714, 1813096560, 1333889218, 700359215, 2002688523, 972070810, 776374577},
    '{244, 857269099, 1772516347, 1560031333, 377198689, 1250286794, 347625639, 1246846107, 115597473, 721409529, 1780062069},
    '{112, 496627171, 1898196697, 299895721, 2123987513, 532972514, 1188892805, 1325819703, 2135574074, 1367990915, 355294580},
    '{164, 1998115579, 1308764907, 85540605, 2013708682, 1749295163, 13950112, 594118444, 735651329, 1579828076, 1823764388},
    '{163, 1674574223, 1641192773, 99654522, 632473956, 1869658600, 1541894688, 1418684196, 1598834793, 277015809, 1457422373},
    '{228, 1282404695, 1505245104, 2093223823, 1648528480, 320151729, 83355351, 1307000805, 1473442512, 1317796606, 2036280055},
    '{22, 2003188085, 899716888, 1871148357, 686871878, 2071732659, 823306320, 75320724, 453239415, 1015068373, 1032114000},
    '{159, 20970055, 1634345209, 2106805199, 2037739287, 1323057583, 1229263839, 1033055347, 376751901, 1999095109, 1495198983},
    '{251, 1483848959, 31822524, 376298145, 154584786, 205551479, 1580451345, 1499335838, 974273047, 433195029, 1789433765},
    '{126, 1581152784, 464912493, 696702010, 2107193264, 1682514016, 220706020, 705519562, 1005951479, 826993455, 1011192223},
    '{175, 1369512941, 329035070, 153233165, 2098761922, 249288194, 2076360433, 1046600320, 1481033675, 1884296552, 351316373},
    '{95, 1568564000, 626777195, 2113275844, 1907172835, 397181129, 1643001689, 1793053262, 1634456268, 953509426, 639062446}
};


`endif
