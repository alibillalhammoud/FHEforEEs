// ================================================================
//  Test-bench :  tb_fastBConvEx_BBa_to_q
//                - ONE deterministic test only
//                - Uses the user-supplied stimulus / answer
// ================================================================
`timescale 1ns/1ps
`include "types.svh"

module tb_fastBConvEx_BBa_to_q;
// ----------------------------------------------------------------
//  DUT I/O
// ----------------------------------------------------------------
logic clk   = 0;
logic reset = 0;
logic in_valid;
logic out_valid;

rns_residue_t input_RNSpoly  [`N_SLOTS][`BBa_BASIS_LEN];   // B‖Ba residues
rns_residue_t output_RNSpoly [`N_SLOTS][`q_BASIS_LEN];     // q residues out

localparam int QLEN     = `q_BASIS_LEN;      // number of q primes
localparam int BBALEN   = `BBa_BASIS_LEN;    // number of B‖Ba primes (input)
// ----------------------------------------------------------------
//  CLOCK
// ----------------------------------------------------------------
always #5 clk = ~clk;

// ----------------------------------------------------------------
//  DUT
// ----------------------------------------------------------------
fastBConvEx_BBa_to_q DUT (
    .clk            (clk),
    .reset          (reset),
    .in_valid       (in_valid),
    .input_RNSpoly  (input_RNSpoly),
    .out_valid      (out_valid),
    .output_RNSpoly (output_RNSpoly)
);

// ----------------------------------------------------------------
//  USER-SUPPLIED TEST VECTORS
// ----------------------------------------------------------------
localparam int NUM_TRIALS = 1;  //  one run only

// test stimulus here
const rns_residue_t KNOWN_IN [`N_SLOTS][`BBa_BASIS_LEN] = '{
    '{2406575, 313906966, 605474624, 934239537, 1589668363, 1567356734, 1471776138, 364225185, 1613769651, 1153893135, 1856411822},
    '{81001096, 511913739, 1130195616, 935905454, 1510787025, 1859042182, 520698806, 141283181, 957394802, 1041317308, 273885315},
    '{2055992580, 1531891891, 1090933461, 572525100, 1245624002, 287953027, 1925629873, 1565019550, 1660605871, 516066792, 1970769398},
    '{680468203, 1402207188, 847597246, 956089897, 1994455403, 402658697, 1729960384, 1444148079, 1247481335, 104546859, 911579519},
    '{1981331186, 270691168, 578111836, 1485776934, 523322228, 1672899391, 581071596, 209906933, 1937820572, 1722258337, 656554988},
    '{1507789192, 1057874066, 1239533268, 1520038621, 618026960, 637922026, 366521069, 1066877968, 154029783, 266603930, 1749384995},
    '{939961214, 1362239244, 258100131, 635551601, 33265343, 1987051861, 1182272113, 963446960, 1728519845, 592150413, 1185632388},
    '{1459793209, 1114861983, 1708067667, 233711142, 1053016725, 1253721065, 1355798783, 45355269, 708739769, 130643320, 396704188},
    '{1235861497, 1141593479, 1040232804, 1310947662, 1551004462, 744998938, 655539971, 802686368, 326224097, 1070548522, 315525028},
    '{719126444, 1986038605, 1624781605, 1205748015, 578864915, 792759487, 1887702220, 1954252474, 842445442, 2041960974, 1171648770},
    '{993668077, 1208123452, 1870638289, 1437634358, 1217623833, 1817907176, 364254771, 2034380733, 1861736132, 1836298811, 1008315771},
    '{531244676, 176969436, 499291796, 919046049, 363811625, 1243783645, 2093180313, 113600263, 1858652316, 1521120752, 766368520},
    '{512137188, 262417205, 753660508, 996624964, 1438329733, 1707058579, 1561088649, 1973453196, 1026946607, 1195063626, 897700266},
    '{1492782280, 1877260613, 725974715, 2114713929, 1886993401, 1006122773, 64064158, 4562261, 389883655, 1452813470, 140368152},
    '{973137646, 448824411, 1273111477, 1073719071, 124623805, 222994203, 676132011, 147163343, 983114351, 1168296970, 1424746320},
    '{1760891879, 489222995, 1161239651, 611599488, 1369000515, 1880566775, 407302070, 1765713593, 1850035282, 1671526585, 650239463},
    '{99592340, 402659615, 1136250757, 153344595, 539961838, 1017773168, 1351528001, 1903210076, 1127800961, 942725257, 2144914371},
    '{356720379, 726306145, 841674202, 1513398140, 1675121933, 2051788094, 1636822034, 1504253498, 677505606, 1726797323, 431762233},
    '{1797078652, 965189296, 2101889306, 2036607256, 1629679618, 1516407549, 647705664, 141529315, 343187844, 1134852132, 793334257},
    '{1697693148, 602810806, 347465435, 585980505, 957143300, 618156830, 727220297, 1091530320, 90661765, 1315135908, 1392059309},
    '{54406186, 1641040526, 172420453, 20348990, 658270238, 380429789, 767586555, 1925354464, 982583157, 783985997, 782395249},
    '{1360751317, 1221793502, 1655693209, 2032112247, 199413, 1102406212, 2074409899, 1391658613, 1232458906, 1413409323, 1984506769},
    '{1015913994, 194203877, 996827189, 1295829275, 2142890934, 1609431404, 1662833724, 24006374, 1029637171, 1162709024, 1076173463},
    '{414133899, 1054077184, 1522311628, 1266050552, 340419067, 92322600, 1952973300, 769560695, 1233956586, 696948476, 1665236991},
    '{1905660568, 108391766, 686072115, 1169578648, 1369767692, 479475575, 1276715384, 1639168422, 197997224, 2122651339, 2106704340},
    '{2146204958, 1893340932, 2033795022, 854911643, 600729427, 1915012376, 475674864, 1944663921, 158512527, 1748072582, 1858882740},
    '{1256330565, 1363158609, 550996612, 965644187, 655911434, 1442701579, 397793942, 804160830, 2023525790, 1485967739, 1986138205},
    '{790536360, 576932890, 408926549, 608054726, 1037418890, 1035668867, 473407492, 1999421932, 402191142, 64965890, 2017865625},
    '{1066811454, 487286723, 1473468771, 91359911, 1741399031, 2091868701, 1989685199, 834080369, 1295874215, 867456099, 1689179528},
    '{1095444225, 1689395509, 454423238, 756358769, 1761802148, 1556338264, 256421482, 752261882, 1563366245, 587761475, 329435887},
    '{704614972, 628351179, 2123456575, 689287272, 1413576382, 1256201973, 1575448078, 413991834, 579738227, 690582911, 1788497851},
    '{1263759218, 1224427145, 497561573, 2041789324, 525661179, 37790758, 1074328797, 1471993313, 1289280764, 1781870380, 1674283996},
    '{734086029, 1496252073, 1545358428, 517601706, 590606257, 1582342532, 2068120328, 169232049, 1451417623, 1918733375, 169362086},
    '{440875221, 211096, 1975290762, 1864165673, 2132420018, 1997881216, 207978271, 297358748, 223630192, 1296401166, 1132842309},
    '{690969991, 425860733, 613422242, 1169018016, 631200332, 1628298016, 471598227, 1590758801, 1642195566, 71755622, 1598666286},
    '{1064509008, 1171851795, 1664557051, 944936064, 532990375, 1362573797, 1041741186, 1822302322, 1031694695, 907367624, 541551278},
    '{399265170, 644856550, 774293876, 1156413635, 1832643562, 66869645, 1810055000, 705985050, 922869234, 482276845, 198385014},
    '{1597192379, 1793492906, 394564745, 1567243632, 1661645748, 854528972, 1307780663, 1171051708, 1279202903, 939443532, 1519436909},
    '{1287479889, 592383651, 757140919, 986077766, 197728418, 1496347989, 1076023385, 310639074, 1944694510, 1841349452, 1781596949},
    '{877293530, 680735415, 1276096439, 1320432424, 682780658, 245032395, 364988159, 393689510, 1414584694, 106383080, 212476702},
    '{76890534, 1463999637, 1682399220, 312822740, 700779533, 1066818239, 1049517706, 1615351145, 1685240303, 335888525, 2080584363},
    '{1276474204, 281092366, 882130565, 1646368213, 1079802398, 530530517, 218465760, 1825414618, 1328024520, 596714516, 1589355981},
    '{1904784871, 2018720024, 826138003, 897162357, 296692050, 624870, 1522206850, 1573945787, 942611545, 699724978, 1480432030},
    '{172168037, 956953317, 1141769605, 124628910, 81326518, 1744788010, 176857354, 702079915, 1192436350, 1420610320, 1013178392},
    '{795428645, 165369361, 1413723967, 317211378, 126869386, 2139089952, 1910725768, 1183584878, 951374247, 212440062, 991754962},
    '{550123113, 1176413791, 943939508, 944683965, 1098339517, 1155793733, 29380478, 1292246679, 1359073312, 1420581464, 115591543},
    '{1097670016, 920110368, 992106981, 392351802, 1741179579, 1504664780, 1083176042, 1607075061, 72701877, 490662662, 375538199},
    '{853297895, 1549249585, 676457627, 1848545344, 386240396, 709855208, 1066061302, 540213286, 2048147107, 1956987137, 927762976},
    '{1323850257, 164774676, 1678604188, 1953881943, 2062196185, 589043076, 1984699685, 524787334, 1956415317, 917888968, 225000876},
    '{727123941, 1010281021, 1547777933, 882506301, 831072733, 103561200, 1934965260, 2096307526, 682153045, 790133528, 1296402548},
    '{1189060403, 998859921, 1777087363, 1599721371, 1517257180, 1791045272, 187718463, 529070739, 1367756034, 735762285, 1164915924},
    '{1642288113, 2149147, 1194360260, 1593755617, 1287594959, 1327956309, 2142396084, 1142970209, 1468627592, 1166401127, 1005490367},
    '{1883487776, 1721982432, 1449901647, 35967890, 167599815, 2042122320, 1994596462, 1576198708, 808116175, 494991200, 1327915565},
    '{1737756517, 75181361, 250878390, 330465822, 2025578758, 1376875783, 388786945, 1658435564, 1633453352, 304563362, 792004994},
    '{1121753646, 1955676666, 2091500489, 236897374, 394681111, 778270610, 1698553150, 1962482671, 506902708, 714000722, 1942692519},
    '{1046961526, 1032807288, 1201942487, 1456638309, 48840388, 372821246, 686716535, 55738262, 2059014790, 1649686815, 431303318},
    '{856024551, 1126229164, 1158287201, 1340354664, 1493953049, 933558923, 1331379471, 1843382751, 2064308379, 2010055463, 1884754857},
    '{569350354, 338377234, 902771092, 267012725, 912847616, 1341904049, 1742999534, 791530456, 266951401, 23151614, 780811672},
    '{445401295, 698297736, 22414416, 1537993602, 731951509, 212997683, 1649163198, 1338983511, 6556059, 609123505, 1419375288},
    '{454542236, 1841160733, 1625951161, 106803849, 1207382414, 1346454852, 1769967665, 1285718905, 60631945, 1661393899, 994437922},
    '{666346933, 489194288, 879451083, 709680126, 2144914019, 1470930075, 1604786121, 1706382111, 1524219264, 1988380883, 1002808500},
    '{1171553528, 1012450913, 438759822, 976368811, 1731737561, 1750967259, 301582012, 1659309318, 1091393147, 60892554, 984982174},
    '{1495411137, 1638380283, 866160050, 790454697, 1753231758, 960718445, 1928281240, 1972799288, 1951001614, 1453127537, 966844749},
    '{1737016703, 598355960, 606607430, 388968163, 1080018074, 238100719, 36803152, 1026589462, 1393076867, 698860141, 1205040083}
};

const rns_residue_t KNOWN_OUT [`N_SLOTS][`q_BASIS_LEN ] = '{
    '{158, 1801396337, 771080194, 1545482434, 1534409644, 1208356101, 1997810206, 414016370, 1837972434, 1246544663, 865006849},
    '{214, 609480513, 722867419, 1413388221, 1522910038, 789514314, 1203772624, 1661722859, 760917651, 1351751619, 589804970},
    '{22, 1253063869, 1391541022, 748315333, 1649333093, 1924359522, 75902126, 367795152, 1540106940, 1553122456, 895914698},
    '{152, 2000434716, 2011511581, 145341502, 1149729491, 443369048, 100845914, 656334509, 608597249, 1884688561, 2089648351},
    '{230, 2144541702, 2075390131, 405289508, 1566418674, 559549721, 380033446, 1043498005, 1123508056, 2018651604, 1355728670},
    '{212, 1677054203, 1897028132, 1260191508, 1819201300, 583722244, 701745705, 1141521185, 1735122, 432250306, 52427481},
    '{202, 1858194972, 404906410, 186386396, 655073713, 462606061, 1622085330, 1648288969, 1578119023, 398543986, 1976101283},
    '{134, 924217006, 498678017, 151099641, 2043316678, 1700369347, 1419186445, 801365078, 707258900, 1367676179, 1819571956},
    '{199, 116849431, 241103215, 1142800802, 1979071411, 329692928, 72678755, 82481210, 1473772782, 994266700, 320582811},
    '{87, 1213855270, 963192960, 1021134861, 126355880, 208640153, 1951028120, 948786284, 994077235, 1596287466, 214431563},
    '{47, 619398504, 1444987741, 618184725, 1407899840, 1617736779, 1767888569, 824321124, 1406188529, 1151357252, 995453260},
    '{80, 189326378, 274067817, 1610693797, 1530753322, 1334737636, 2143251596, 1129915921, 955464511, 856842171, 1433592267},
    '{192, 115928855, 1305801653, 126122593, 1984399284, 2136675677, 1259369365, 115960391, 1525135389, 640475483, 1441263522},
    '{209, 30716288, 903505795, 2143888487, 1678342436, 427400267, 135650988, 1658953739, 596066332, 2093172133, 1504624300},
    '{91, 197105913, 1407846172, 2096109748, 1831233930, 767550643, 2019405013, 1823108986, 543603311, 1560696287, 1101922330},
    '{137, 575800371, 863707673, 387485420, 718699122, 1867426900, 1806123924, 398333997, 1385160706, 1528953171, 890394004},
    '{27, 1721613664, 1265017699, 1577603838, 341769223, 908151536, 1696092013, 95410762, 1988723855, 768096938, 136253847},
    '{128, 1641060792, 111535544, 966644686, 1485718645, 1308398528, 2025713005, 756470905, 190171630, 402554121, 1354868192},
    '{37, 292087364, 122652427, 764407335, 1225851744, 1833407878, 1145178764, 1787282124, 1395632859, 1666944916, 1413646642},
    '{223, 311482435, 55223871, 1132294007, 872954559, 963561611, 645731369, 1653343971, 506343028, 118178695, 1390687547},
    '{60, 617058589, 1753332016, 1165613387, 533351539, 1820292411, 2021621146, 540154887, 498055378, 536055491, 482518146},
    '{183, 1997261724, 762031393, 1446043103, 795679453, 67225453, 1115426426, 498403647, 888362128, 1532621427, 1458534471},
    '{193, 402910588, 1465683659, 1247326843, 2134297682, 390455062, 1304105150, 1781585723, 1735051744, 561538982, 296227189},
    '{239, 2003485789, 1845605540, 577868776, 336652826, 394557723, 1574337103, 1961626260, 2089727793, 1051929917, 1400360844},
    '{55, 221134128, 955390720, 1132368144, 1173180839, 1458333344, 954294901, 557036859, 2115164745, 1983792286, 123016169},
    '{30, 1386746641, 1335526754, 950421705, 602345192, 752812172, 128946916, 1193232123, 1899808246, 1887933193, 1409526560},
    '{241, 1043780466, 847578797, 1303964814, 455721696, 100342289, 1934730061, 123370419, 1059132888, 385943998, 1588078904},
    '{85, 1303166692, 393147312, 566898218, 702283574, 1868992300, 245029595, 1024497426, 570417274, 1821432966, 231691757},
    '{44, 700917930, 859089615, 2049229424, 2061297855, 1971226300, 751506102, 1705141657, 2131048474, 1218447018, 608686242},
    '{237, 1862133786, 1036391050, 1855291657, 1156636861, 1745498165, 1920691979, 430507648, 974571625, 323475878, 1636889060},
    '{253, 2015055566, 1857652332, 1714673096, 1630710979, 716443577, 444735163, 750022632, 439239608, 1170533342, 1393903665},
    '{103, 1470627387, 105414309, 1204875268, 1627894244, 1682718118, 2118395920, 601864015, 107809099, 1024055309, 538944420},
    '{205, 389526391, 767297735, 2133167035, 2052513320, 545086098, 1462428058, 720688122, 1348990143, 87660997, 191374085},
    '{126, 1104566358, 1853491678, 1644961877, 1693302834, 2027966286, 171539455, 902926787, 1692012824, 1002430574, 108734014},
    '{253, 2146905725, 1976014662, 439795418, 1371243517, 1706485710, 980519577, 1883616662, 11887144, 1569415834, 1545188894},
    '{230, 1448990006, 301223854, 1670525462, 1549897681, 764220675, 1692620784, 1776542014, 1420991268, 1045544343, 258651919},
    '{167, 1415823220, 1171314222, 568379186, 1243515384, 1984897333, 486859124, 1502576021, 767284067, 1260932241, 958250409},
    '{34, 1904635914, 2078243115, 1999510873, 2026157157, 378901098, 38207575, 162912908, 982499901, 31548800, 419028592},
    '{149, 170762404, 95215766, 608831440, 1917924280, 909053913, 2090585190, 2053131771, 1301788880, 654717821, 84751483},
    '{118, 1804546386, 204586843, 161228441, 1150884585, 2013435374, 1506243889, 112026913, 1464663341, 1597035310, 1975756930},
    '{42, 93184485, 1800513439, 207225707, 1358240790, 1750089657, 1588644679, 1788503073, 1639771590, 1865438283, 1439225757},
    '{9, 1202563950, 893945767, 1607297058, 1354676769, 190537601, 401453242, 1716216147, 1239399530, 1032772819, 1572771833},
    '{218, 711737088, 310049076, 1499327940, 2100764522, 1556288262, 130741760, 652332428, 395627464, 990540216, 777903151},
    '{4, 28956712, 1826064697, 1269978679, 961265842, 1477047224, 1799274657, 1566364137, 194928113, 592821815, 2134909736},
    '{207, 1161637796, 547561824, 1138257451, 2034390903, 1642658467, 976063638, 1256471042, 108710816, 239982289, 632608984},
    '{65, 1037658993, 1455334569, 653284961, 1723592142, 1295944025, 1871635865, 357089516, 1313109111, 298369002, 432738018},
    '{58, 276987747, 1822728999, 1412869425, 1254383419, 878122169, 1000302496, 962329306, 718919697, 356678555, 434814004},
    '{155, 313366688, 1338392354, 725318873, 488045733, 1036207313, 1985581360, 41064856, 487185765, 402883747, 2085083490},
    '{208, 197470081, 1652161501, 1568782751, 245772867, 1395996992, 701114206, 1036673856, 788221428, 378554379, 1722989319},
    '{82, 795968331, 1385102178, 1492702467, 411407149, 1465398324, 1994328464, 1197423838, 1058462584, 1626028574, 1914681308},
    '{211, 1366114, 1043855037, 670333125, 1198628788, 1285567930, 2098576741, 1850785061, 685521850, 346864839, 1357249972},
    '{64, 1280752672, 497276370, 1563371972, 1975234218, 263011793, 636260153, 1099600829, 1805754923, 1145337591, 1037881926},
    '{72, 1978056554, 138183431, 2136438202, 544797235, 1145809227, 143343672, 1768436228, 1763843905, 1125580866, 1432344677},
    '{239, 36559424, 1068305945, 291205652, 1950603649, 1810800871, 12863017, 459252221, 1023501629, 581696926, 2044648128},
    '{65, 830131868, 441235074, 843785352, 672304345, 1548466971, 1701404323, 1346631372, 319034943, 1954077396, 7073732},
    '{226, 632447839, 1084997531, 1649095537, 414106287, 1649923524, 31532308, 725927437, 124455211, 71844703, 1418781788},
    '{195, 845394424, 1953615215, 912150056, 426821088, 1744749443, 1798743154, 1396512290, 1373770693, 684046346, 1244813943},
    '{6, 1685871322, 1870169621, 1319915917, 1554012325, 1959965337, 1463540128, 1781629019, 1533809718, 1500726479, 1208865636},
    '{136, 1698647832, 330866251, 754632812, 2038023307, 814813097, 1072222957, 889400428, 1696919904, 2055134257, 1963350687},
    '{104, 1480075337, 583237565, 1597096057, 1605215835, 1150390998, 125693025, 597560394, 2142732665, 968489025, 1544833141},
    '{77, 168947452, 251594094, 1577034622, 1279223584, 1522438008, 1130549699, 878140950, 1109346268, 1918644444, 1597702600},
    '{252, 2110522965, 1059776876, 113313473, 1925142556, 32071784, 816480111, 545969148, 518243365, 1452923143, 102471743},
    '{110, 82806304, 1800884278, 1287556023, 1502521424, 773486774, 1268138829, 448977532, 1327512067, 856409846, 1457182071},
    '{0, 1821404230, 2008770391, 1214484748, 1190232239, 233720945, 1124115358, 2024202829, 117897968, 1815038935, 1489867147}
};


// ----------------------------------------------------------------
//  TEST PROGRAM
// ----------------------------------------------------------------
rns_residue_t golden_answer [`N_SLOTS][`q_BASIS_LEN];
bit           mismatch;
int unsigned  pass_cnt = 0;
int unsigned  fail_cnt = 0;
logic DEBUG_MODE = 0;

initial begin
   // ------------- reset sequence -------------
   @(posedge clk);
   @(negedge clk);
   reset    = 1'b1;
   in_valid = 1'b0;
   @(negedge clk);
   reset    = 1'b0;

   // *************************************************************
   //  ONLY ONE TRIAL – load the static vectors
   // *************************************************************
   for (int k = 0; k < `N_SLOTS; k++) begin
      // copy the whole B‖Ba basis
      for (int j = 0; j < BBALEN; j++) begin
         input_RNSpoly[k][j]  = KNOWN_IN [k][j];
      end
      // copy expected q-basis answer
      for (int j = 0; j < QLEN; j++) begin
         golden_answer[k][j]  = KNOWN_OUT[k][j];
      end
   end

   // -------------- Drive DUT -----------------
   @(negedge clk);
   in_valid = 1'b1;
   @(negedge clk);
   in_valid = 1'b0;

   if (DEBUG_MODE) begin
      // Display [1][1] and [1][2] for input_RNSpoly and output_RNSpoly
      $display("[%0t] input_RNSpoly[1][1]=%0d  input_RNSpoly[1][2]=%0d", $time, DUT.input_RNSpoly[1][1], DUT.input_RNSpoly[1][2]);
      //$monitor("[%0t] output_RNSpoly[1][1]=%0d  output_RNSpoly[1][2]=%0d", $time, DUT.output_RNSpoly[1][1], DUT.output_RNSpoly[1][2]);
      //$monitor("[%0t] temp[1]=%0d gamma[1]=%0d", $time, DUT.temp[1], DUT.gamma_centered[1]);
      //$monitor("[%0t] xB_to_q[1][1]=%0d", $time, DUT.xB_in_q[1][1]);
      //$monitor("[%0t] rr_tmpvar1[1][1]=%0d", $time, DUT.rr_tmpvar1[1][1]);
      $monitor("[%0t] rr_tmpvar2[1][1]=%0d , rr_tmpvar3[1][1]=%0d", $time, DUT.rr_tmpvar2[1][1], DUT.rr_tmpvar3_mod[1][1]);
      //$monitor("[%0t] rr_tmpvar3[1][1]=%0d", $time, DUT.rr_tmpvar3_mod[1][1]);
      // If you want to look inside the DUT at intermediate signals, try (if public in your module):
      //$monitor("[%0t] DUT.xB_RNSpoly[1][1]=%0d  DUT.xB_RNSpoly[1][2]=%0d", $time, DUT.xB_RNSpoly[1][1], DUT.xB_RNSpoly[1][2]);
      //$monitor("[%0t] DUT.xB_in_q[1][1]=%0d  DUT.xB_in_q[1][2]=%0d", $time, DUT.xB_in_q[1][1], DUT.xB_in_q[1][2]);
   end
   //$display("[%0t] xB_RNSpoly[1][1]=%0d  signed_xBa_RNSpoly[1][0]=%0d", $time, DUT.xB_RNSpoly[1][1], DUT.signed_xBa_RNSpoly[1][0]);


   // -------------- Wait for result -----------
   while (!out_valid) @(posedge clk);
   //$display("[%0t] rr_tmpvar2[1][1] mod qbasis[1] = %0d", $time, DUT.rr_tmpvar2[1][1] % q_BASIS[1]);

   // -------------- Compare -------------------
   mismatch = 0;
   for (int k = 0; k < `N_SLOTS; k++) begin
      for (int j = 0; j < QLEN; j++) begin
         if (output_RNSpoly[k][j] !== golden_answer[k][j]) begin
            $display("[%0t]  SLOT %0d  RES %0d  MISMATCH  DUT=%0d  GOLD=%0d", $time, k, j, output_RNSpoly[k][j], golden_answer[k][j]);
            mismatch = 1;
         end
      end
   end
   //$display("[%0t] output_RNSpoly[1][1]=%0d  output_RNSpoly[1][2]=%0d", $time, DUT.output_RNSpoly[1][1], DUT.output_RNSpoly[1][2]);

   if (mismatch) fail_cnt++; else pass_cnt++;

   // -------------- Summary -------------------
   $display("\n==================================================");
   $display("fastBConvEx deterministic test finished");
   $display("      Passed : %0d", pass_cnt);
   $display("      Failed : %0d", fail_cnt);
   $display("==================================================\n");
   $finish;
end

endmodule